// Generator : SpinalHDL v1.6.4    git head : 598c18959149eb18e5eee5b0aa3eef01ecaa41a1
// Component : PoseidonTopLevel

`timescale 1ns/1ps 

module PoseidonTopLevel (
  input               io_input_valid,
  output              io_input_ready,
  input               io_input_last,
  input      [254:0]  io_input_payload,
  output              io_output_valid,
  input               io_output_ready,
  output              io_output_last,
  output     [254:0]  io_output_payload,
  input               clk,
  input               resetn
);
import "DPI-C" function void c_py_gen_packet(output bit[255:0] pkt);

  reg                 poseidonLoop_1_io_output_ready;
  wire                aXI4StreamReceiver_1_io_input_ready;
  wire                aXI4StreamReceiver_1_io_output_valid;
  wire                aXI4StreamReceiver_1_io_output_payload_isFull;
  wire       [2:0]    aXI4StreamReceiver_1_io_output_payload_fullRound;
  wire       [5:0]    aXI4StreamReceiver_1_io_output_payload_partialRound;
  wire       [3:0]    aXI4StreamReceiver_1_io_output_payload_stateSize;
  wire       [7:0]    aXI4StreamReceiver_1_io_output_payload_stateID;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_0;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_1;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_2;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_3;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_4;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_5;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_6;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_7;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_8;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_9;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_10;
  wire       [254:0]  aXI4StreamReceiver_1_io_output_payload_stateElements_11;
  wire                poseidonLoop_1_io_input_ready;
  wire                poseidonLoop_1_io_output_valid;
  wire       [7:0]    poseidonLoop_1_io_output_payload_stateID;
  wire       [254:0]  poseidonLoop_1_io_output_payload_stateElement;
  wire                aXI4StreamTransmitter_1_io_input_ready;
  wire                aXI4StreamTransmitter_1_io_output_valid;
  wire                aXI4StreamTransmitter_1_io_output_last;
  wire       [254:0]  aXI4StreamTransmitter_1_io_output_payload;
  wire                poseidonLoop_1_io_output_m2sPipe_valid;
  wire                poseidonLoop_1_io_output_m2sPipe_ready;
  wire       [7:0]    poseidonLoop_1_io_output_m2sPipe_payload_stateID;
  wire       [254:0]  poseidonLoop_1_io_output_m2sPipe_payload_stateElement;
  reg                 poseidonLoop_1_io_output_rValid;
  reg        [7:0]    poseidonLoop_1_io_output_rData_stateID;
  reg        [254:0]  poseidonLoop_1_io_output_rData_stateElement;
  wire                when_Stream_l342;

  AXI4StreamReceiver aXI4StreamReceiver_1 (
    .io_input_valid                        (io_input_valid                                                  ), //i
    .io_input_ready                        (aXI4StreamReceiver_1_io_input_ready                             ), //o
    .io_input_last                         (io_input_last                                                   ), //i
    .io_input_payload                      (io_input_payload[254:0]                                         ), //i
    .io_output_valid                       (aXI4StreamReceiver_1_io_output_valid                            ), //o
    .io_output_ready                       (poseidonLoop_1_io_input_ready                                   ), //i
    .io_output_payload_isFull              (aXI4StreamReceiver_1_io_output_payload_isFull                   ), //o
    .io_output_payload_fullRound           (aXI4StreamReceiver_1_io_output_payload_fullRound[2:0]           ), //o
    .io_output_payload_partialRound        (aXI4StreamReceiver_1_io_output_payload_partialRound[5:0]        ), //o
    .io_output_payload_stateSize           (aXI4StreamReceiver_1_io_output_payload_stateSize[3:0]           ), //o
    .io_output_payload_stateID             (aXI4StreamReceiver_1_io_output_payload_stateID[7:0]             ), //o
    .io_output_payload_stateElements_0     (aXI4StreamReceiver_1_io_output_payload_stateElements_0[254:0]   ), //o
    .io_output_payload_stateElements_1     (aXI4StreamReceiver_1_io_output_payload_stateElements_1[254:0]   ), //o
    .io_output_payload_stateElements_2     (aXI4StreamReceiver_1_io_output_payload_stateElements_2[254:0]   ), //o
    .io_output_payload_stateElements_3     (aXI4StreamReceiver_1_io_output_payload_stateElements_3[254:0]   ), //o
    .io_output_payload_stateElements_4     (aXI4StreamReceiver_1_io_output_payload_stateElements_4[254:0]   ), //o
    .io_output_payload_stateElements_5     (aXI4StreamReceiver_1_io_output_payload_stateElements_5[254:0]   ), //o
    .io_output_payload_stateElements_6     (aXI4StreamReceiver_1_io_output_payload_stateElements_6[254:0]   ), //o
    .io_output_payload_stateElements_7     (aXI4StreamReceiver_1_io_output_payload_stateElements_7[254:0]   ), //o
    .io_output_payload_stateElements_8     (aXI4StreamReceiver_1_io_output_payload_stateElements_8[254:0]   ), //o
    .io_output_payload_stateElements_9     (aXI4StreamReceiver_1_io_output_payload_stateElements_9[254:0]   ), //o
    .io_output_payload_stateElements_10    (aXI4StreamReceiver_1_io_output_payload_stateElements_10[254:0]  ), //o
    .io_output_payload_stateElements_11    (aXI4StreamReceiver_1_io_output_payload_stateElements_11[254:0]  ), //o
    .clk                                   (clk                                                             ), //i
    .resetn                                (resetn                                                          )  //i
  );
  PoseidonLoop poseidonLoop_1 (
    .io_input_valid                       (aXI4StreamReceiver_1_io_output_valid                            ), //i
    .io_input_ready                       (poseidonLoop_1_io_input_ready                                   ), //o
    .io_input_payload_isFull              (aXI4StreamReceiver_1_io_output_payload_isFull                   ), //i
    .io_input_payload_fullRound           (aXI4StreamReceiver_1_io_output_payload_fullRound[2:0]           ), //i
    .io_input_payload_partialRound        (aXI4StreamReceiver_1_io_output_payload_partialRound[5:0]        ), //i
    .io_input_payload_stateSize           (aXI4StreamReceiver_1_io_output_payload_stateSize[3:0]           ), //i
    .io_input_payload_stateID             (aXI4StreamReceiver_1_io_output_payload_stateID[7:0]             ), //i
    .io_input_payload_stateElements_0     (aXI4StreamReceiver_1_io_output_payload_stateElements_0[254:0]   ), //i
    .io_input_payload_stateElements_1     (aXI4StreamReceiver_1_io_output_payload_stateElements_1[254:0]   ), //i
    .io_input_payload_stateElements_2     (aXI4StreamReceiver_1_io_output_payload_stateElements_2[254:0]   ), //i
    .io_input_payload_stateElements_3     (aXI4StreamReceiver_1_io_output_payload_stateElements_3[254:0]   ), //i
    .io_input_payload_stateElements_4     (aXI4StreamReceiver_1_io_output_payload_stateElements_4[254:0]   ), //i
    .io_input_payload_stateElements_5     (aXI4StreamReceiver_1_io_output_payload_stateElements_5[254:0]   ), //i
    .io_input_payload_stateElements_6     (aXI4StreamReceiver_1_io_output_payload_stateElements_6[254:0]   ), //i
    .io_input_payload_stateElements_7     (aXI4StreamReceiver_1_io_output_payload_stateElements_7[254:0]   ), //i
    .io_input_payload_stateElements_8     (aXI4StreamReceiver_1_io_output_payload_stateElements_8[254:0]   ), //i
    .io_input_payload_stateElements_9     (aXI4StreamReceiver_1_io_output_payload_stateElements_9[254:0]   ), //i
    .io_input_payload_stateElements_10    (aXI4StreamReceiver_1_io_output_payload_stateElements_10[254:0]  ), //i
    .io_input_payload_stateElements_11    (aXI4StreamReceiver_1_io_output_payload_stateElements_11[254:0]  ), //i
    .io_output_valid                      (poseidonLoop_1_io_output_valid                                  ), //o
    .io_output_ready                      (poseidonLoop_1_io_output_ready                                  ), //i
    .io_output_payload_stateID            (poseidonLoop_1_io_output_payload_stateID[7:0]                   ), //o
    .io_output_payload_stateElement       (poseidonLoop_1_io_output_payload_stateElement[254:0]            ), //o
    .clk                                  (clk                                                             ), //i
    .resetn                               (resetn                                                          )  //i
  );
  AXI4StreamTransmitter aXI4StreamTransmitter_1 (
    .io_input_valid                   (poseidonLoop_1_io_output_m2sPipe_valid                        ), //i
    .io_input_ready                   (aXI4StreamTransmitter_1_io_input_ready                        ), //o
    .io_input_payload_stateID         (poseidonLoop_1_io_output_m2sPipe_payload_stateID[7:0]         ), //i
    .io_input_payload_stateElement    (poseidonLoop_1_io_output_m2sPipe_payload_stateElement[254:0]  ), //i
    .io_output_valid                  (aXI4StreamTransmitter_1_io_output_valid                       ), //o
    .io_output_ready                  (io_output_ready                                               ), //i
    .io_output_last                   (aXI4StreamTransmitter_1_io_output_last                        ), //o
    .io_output_payload                (aXI4StreamTransmitter_1_io_output_payload[254:0]              ), //o
    .clk                              (clk                                                           ), //i
    .resetn                           (resetn                                                        )  //i
  );
  assign io_input_ready = aXI4StreamReceiver_1_io_input_ready;
  always @(*) begin
    poseidonLoop_1_io_output_ready = poseidonLoop_1_io_output_m2sPipe_ready;
    if(when_Stream_l342) begin
      poseidonLoop_1_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! poseidonLoop_1_io_output_m2sPipe_valid);
  assign poseidonLoop_1_io_output_m2sPipe_valid = poseidonLoop_1_io_output_rValid;
  assign poseidonLoop_1_io_output_m2sPipe_payload_stateID = poseidonLoop_1_io_output_rData_stateID;
  assign poseidonLoop_1_io_output_m2sPipe_payload_stateElement = poseidonLoop_1_io_output_rData_stateElement;
  assign poseidonLoop_1_io_output_m2sPipe_ready = aXI4StreamTransmitter_1_io_input_ready;
  assign io_output_valid = aXI4StreamTransmitter_1_io_output_valid;
  assign io_output_last = aXI4StreamTransmitter_1_io_output_last;
  assign io_output_payload = aXI4StreamTransmitter_1_io_output_payload;
  always @(posedge clk) begin
    if(!resetn) begin
      poseidonLoop_1_io_output_rValid <= 1'b0;
    end else begin
      if(poseidonLoop_1_io_output_ready) begin
        poseidonLoop_1_io_output_rValid <= poseidonLoop_1_io_output_valid;
      end
    end
  end

  always @(posedge clk) begin
    if(poseidonLoop_1_io_output_ready) begin
      poseidonLoop_1_io_output_rData_stateID <= poseidonLoop_1_io_output_payload_stateID;
      poseidonLoop_1_io_output_rData_stateElement <= poseidonLoop_1_io_output_payload_stateElement;
    end
  end


endmodule

module AXI4StreamTransmitter (
  input               io_input_valid,
  output              io_input_ready,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElement,
  output              io_output_valid,
  input               io_output_ready,
  output              io_output_last,
  output     [254:0]  io_output_payload,
  input               clk,
  input               resetn
);

  reg                 streamArbiter_2_io_output_ready;
  wire       [0:0]    streamDemux_2_io_select;
  wire                streamDemux_2_io_outputs_0_fifo_io_pop_ready;
  wire                streamArbiter_2_io_inputs_0_ready;
  wire                streamArbiter_2_io_inputs_1_ready;
  wire                streamArbiter_2_io_output_valid;
  wire       [7:0]    streamArbiter_2_io_output_payload_stateID;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElement;
  wire       [0:0]    streamArbiter_2_io_chosen;
  wire       [1:0]    streamArbiter_2_io_chosenOH;
  wire                streamDemux_2_io_input_ready;
  wire                streamDemux_2_io_outputs_0_valid;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_stateID;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElement;
  wire                streamDemux_2_io_outputs_1_valid;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_stateID;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElement;
  wire                streamDemux_2_io_outputs_0_fifo_io_push_ready;
  wire                streamDemux_2_io_outputs_0_fifo_io_pop_valid;
  wire       [7:0]    streamDemux_2_io_outputs_0_fifo_io_pop_payload_stateID;
  wire       [254:0]  streamDemux_2_io_outputs_0_fifo_io_pop_payload_stateElement;
  wire       [3:0]    streamDemux_2_io_outputs_0_fifo_io_occupancy;
  wire       [3:0]    streamDemux_2_io_outputs_0_fifo_io_availability;
  reg        [7:0]    idCounter;
  wire                when_AXI4StreamInterface_l103;
  wire                loopback_valid;
  wire                loopback_ready;
  wire       [7:0]    loopback_payload_stateID;
  wire       [254:0]  loopback_payload_stateElement;
  wire                temp_valid;
  wire                temp_ready;
  wire       [7:0]    temp_payload_stateID;
  wire       [254:0]  temp_payload_stateElement;
  reg                 streamArbiter_2_io_output_rValid;
  reg        [7:0]    streamArbiter_2_io_output_rData_stateID;
  reg        [254:0]  streamArbiter_2_io_output_rData_stateElement;
  wire                when_Stream_l342;
  wire                streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_valid;
  wire                streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_ready;
  wire       [7:0]    streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_payload_stateID;
  wire       [254:0]  streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_payload_stateElement;
  reg                 streamDemux_2_io_outputs_0_fifo_io_pop_rValid;
  reg        [7:0]    streamDemux_2_io_outputs_0_fifo_io_pop_rData_stateID;
  reg        [254:0]  streamDemux_2_io_outputs_0_fifo_io_pop_rData_stateElement;

  StreamArbiter_1 streamArbiter_2 (
    .io_inputs_0_valid                   (io_input_valid                                         ), //i
    .io_inputs_0_ready                   (streamArbiter_2_io_inputs_0_ready                      ), //o
    .io_inputs_0_payload_stateID         (io_input_payload_stateID[7:0]                          ), //i
    .io_inputs_0_payload_stateElement    (io_input_payload_stateElement[254:0]                   ), //i
    .io_inputs_1_valid                   (loopback_valid                                         ), //i
    .io_inputs_1_ready                   (streamArbiter_2_io_inputs_1_ready                      ), //o
    .io_inputs_1_payload_stateID         (loopback_payload_stateID[7:0]                          ), //i
    .io_inputs_1_payload_stateElement    (loopback_payload_stateElement[254:0]                   ), //i
    .io_output_valid                     (streamArbiter_2_io_output_valid                        ), //o
    .io_output_ready                     (streamArbiter_2_io_output_ready                        ), //i
    .io_output_payload_stateID           (streamArbiter_2_io_output_payload_stateID[7:0]         ), //o
    .io_output_payload_stateElement      (streamArbiter_2_io_output_payload_stateElement[254:0]  ), //o
    .io_chosen                           (streamArbiter_2_io_chosen                              ), //o
    .io_chosenOH                         (streamArbiter_2_io_chosenOH[1:0]                       ), //o
    .clk                                 (clk                                                    ), //i
    .resetn                              (resetn                                                 )  //i
  );
  StreamDemux_1 streamDemux_2 (
    .io_select                            (streamDemux_2_io_select                                 ), //i
    .io_input_valid                       (temp_valid                                              ), //i
    .io_input_ready                       (streamDemux_2_io_input_ready                            ), //o
    .io_input_payload_stateID             (temp_payload_stateID[7:0]                               ), //i
    .io_input_payload_stateElement        (temp_payload_stateElement[254:0]                        ), //i
    .io_outputs_0_valid                   (streamDemux_2_io_outputs_0_valid                        ), //o
    .io_outputs_0_ready                   (streamDemux_2_io_outputs_0_fifo_io_push_ready           ), //i
    .io_outputs_0_payload_stateID         (streamDemux_2_io_outputs_0_payload_stateID[7:0]         ), //o
    .io_outputs_0_payload_stateElement    (streamDemux_2_io_outputs_0_payload_stateElement[254:0]  ), //o
    .io_outputs_1_valid                   (streamDemux_2_io_outputs_1_valid                        ), //o
    .io_outputs_1_ready                   (io_output_ready                                         ), //i
    .io_outputs_1_payload_stateID         (streamDemux_2_io_outputs_1_payload_stateID[7:0]         ), //o
    .io_outputs_1_payload_stateElement    (streamDemux_2_io_outputs_1_payload_stateElement[254:0]  )  //o
  );
  StreamFifo_1 streamDemux_2_io_outputs_0_fifo (
    .io_push_valid                   (streamDemux_2_io_outputs_0_valid                                    ), //i
    .io_push_ready                   (streamDemux_2_io_outputs_0_fifo_io_push_ready                       ), //o
    .io_push_payload_stateID         (streamDemux_2_io_outputs_0_payload_stateID[7:0]                     ), //i
    .io_push_payload_stateElement    (streamDemux_2_io_outputs_0_payload_stateElement[254:0]              ), //i
    .io_pop_valid                    (streamDemux_2_io_outputs_0_fifo_io_pop_valid                        ), //o
    .io_pop_ready                    (streamDemux_2_io_outputs_0_fifo_io_pop_ready                        ), //i
    .io_pop_payload_stateID          (streamDemux_2_io_outputs_0_fifo_io_pop_payload_stateID[7:0]         ), //o
    .io_pop_payload_stateElement     (streamDemux_2_io_outputs_0_fifo_io_pop_payload_stateElement[254:0]  ), //o
    .io_flush                        (1'b0                                                                ), //i
    .io_occupancy                    (streamDemux_2_io_outputs_0_fifo_io_occupancy[3:0]                   ), //o
    .io_availability                 (streamDemux_2_io_outputs_0_fifo_io_availability[3:0]                ), //o
    .clk                             (clk                                                                 ), //i
    .resetn                          (resetn                                                              )  //i
  );
  assign when_AXI4StreamInterface_l103 = (io_output_valid && io_output_ready);
  assign io_input_ready = streamArbiter_2_io_inputs_0_ready;
  assign loopback_ready = streamArbiter_2_io_inputs_1_ready;
  always @(*) begin
    streamArbiter_2_io_output_ready = temp_ready;
    if(when_Stream_l342) begin
      streamArbiter_2_io_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! temp_valid);
  assign temp_valid = streamArbiter_2_io_output_rValid;
  assign temp_payload_stateID = streamArbiter_2_io_output_rData_stateID;
  assign temp_payload_stateElement = streamArbiter_2_io_output_rData_stateElement;
  assign temp_ready = streamDemux_2_io_input_ready;
  assign streamDemux_2_io_select = (temp_payload_stateID == idCounter);
  assign io_output_last = 1'b1;
  assign io_output_valid = streamDemux_2_io_outputs_1_valid;
  assign io_output_payload = streamDemux_2_io_outputs_1_payload_stateElement;
  assign streamDemux_2_io_outputs_0_fifo_io_pop_ready = (! streamDemux_2_io_outputs_0_fifo_io_pop_rValid);
  assign streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_valid = (streamDemux_2_io_outputs_0_fifo_io_pop_valid || streamDemux_2_io_outputs_0_fifo_io_pop_rValid);
  assign streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_payload_stateID = (streamDemux_2_io_outputs_0_fifo_io_pop_rValid ? streamDemux_2_io_outputs_0_fifo_io_pop_rData_stateID : streamDemux_2_io_outputs_0_fifo_io_pop_payload_stateID);
  assign streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_payload_stateElement = (streamDemux_2_io_outputs_0_fifo_io_pop_rValid ? streamDemux_2_io_outputs_0_fifo_io_pop_rData_stateElement : streamDemux_2_io_outputs_0_fifo_io_pop_payload_stateElement);
  assign loopback_valid = streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_valid;
  assign streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_ready = loopback_ready;
  assign loopback_payload_stateID = streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_payload_stateID;
  assign loopback_payload_stateElement = streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_payload_stateElement;
  always @(posedge clk) begin
    if(!resetn) begin
      idCounter <= 8'h0;
      streamArbiter_2_io_output_rValid <= 1'b0;
      streamDemux_2_io_outputs_0_fifo_io_pop_rValid <= 1'b0;
    end else begin
      if(when_AXI4StreamInterface_l103) begin
        idCounter <= (idCounter + 8'h01);
      end
      if(streamArbiter_2_io_output_ready) begin
        streamArbiter_2_io_output_rValid <= streamArbiter_2_io_output_valid;
      end
      if(streamDemux_2_io_outputs_0_fifo_io_pop_valid) begin
        streamDemux_2_io_outputs_0_fifo_io_pop_rValid <= 1'b1;
      end
      if(streamDemux_2_io_outputs_0_fifo_io_pop_s2mPipe_ready) begin
        streamDemux_2_io_outputs_0_fifo_io_pop_rValid <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(streamArbiter_2_io_output_ready) begin
      streamArbiter_2_io_output_rData_stateID <= streamArbiter_2_io_output_payload_stateID;
      streamArbiter_2_io_output_rData_stateElement <= streamArbiter_2_io_output_payload_stateElement;
    end
    if(streamDemux_2_io_outputs_0_fifo_io_pop_ready) begin
      streamDemux_2_io_outputs_0_fifo_io_pop_rData_stateID <= streamDemux_2_io_outputs_0_fifo_io_pop_payload_stateID;
      streamDemux_2_io_outputs_0_fifo_io_pop_rData_stateElement <= streamDemux_2_io_outputs_0_fifo_io_pop_payload_stateElement;
    end
  end


endmodule

module PoseidonLoop (
  input               io_input_valid,
  output              io_input_ready,
  input               io_input_payload_isFull,
  input      [2:0]    io_input_payload_fullRound,
  input      [5:0]    io_input_payload_partialRound,
  input      [3:0]    io_input_payload_stateSize,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElements_0,
  input      [254:0]  io_input_payload_stateElements_1,
  input      [254:0]  io_input_payload_stateElements_2,
  input      [254:0]  io_input_payload_stateElements_3,
  input      [254:0]  io_input_payload_stateElements_4,
  input      [254:0]  io_input_payload_stateElements_5,
  input      [254:0]  io_input_payload_stateElements_6,
  input      [254:0]  io_input_payload_stateElements_7,
  input      [254:0]  io_input_payload_stateElements_8,
  input      [254:0]  io_input_payload_stateElements_9,
  input      [254:0]  io_input_payload_stateElements_10,
  input      [254:0]  io_input_payload_stateElements_11,
  output              io_output_valid,
  input               io_output_ready,
  output     [7:0]    io_output_payload_stateID,
  output     [254:0]  io_output_payload_stateElement,
  input               clk,
  input               resetn
);

  wire                demuxInst_io_output0_ready;
  reg                 demuxInst_io_output1_ready;
  wire                streamArbiter_2_io_inputs_0_ready;
  wire                streamArbiter_2_io_inputs_1_ready;
  wire                streamArbiter_2_io_output_valid;
  wire                streamArbiter_2_io_output_payload_isFull;
  wire       [2:0]    streamArbiter_2_io_output_payload_fullRound;
  wire       [5:0]    streamArbiter_2_io_output_payload_partialRound;
  wire       [3:0]    streamArbiter_2_io_output_payload_stateSize;
  wire       [7:0]    streamArbiter_2_io_output_payload_stateID;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_0;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_1;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_2;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_3;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_4;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_5;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_6;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_7;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_8;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_9;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_10;
  wire       [254:0]  streamArbiter_2_io_output_payload_stateElements_11;
  wire       [0:0]    streamArbiter_2_io_chosen;
  wire       [1:0]    streamArbiter_2_io_chosenOH;
  wire                poseidonSerializer_1_io_input_ready;
  wire                poseidonSerializer_1_io_output_valid;
  wire                poseidonSerializer_1_io_output_payload_isFull;
  wire       [2:0]    poseidonSerializer_1_io_output_payload_fullRound;
  wire       [5:0]    poseidonSerializer_1_io_output_payload_partialRound;
  wire       [3:0]    poseidonSerializer_1_io_output_payload_stateIndex;
  wire       [3:0]    poseidonSerializer_1_io_output_payload_stateSize;
  wire       [7:0]    poseidonSerializer_1_io_output_payload_stateID;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_0;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_1;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_2;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_3;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_4;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_5;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_6;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_7;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_8;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_9;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElements_10;
  wire       [254:0]  poseidonSerializer_1_io_output_payload_stateElement;
  wire       [254:0]  preRoundConstantMem_1_io_preConstant;
  wire                preRoundConstStage_adderInst_io_output_valid;
  wire       [254:0]  preRoundConstStage_adderInst_io_output_payload_res;
  wire                poseidonThread_1_io_output_valid;
  wire                poseidonThread_1_io_output_payload_isFull;
  wire       [2:0]    poseidonThread_1_io_output_payload_fullRound;
  wire       [5:0]    poseidonThread_1_io_output_payload_partialRound;
  wire       [3:0]    poseidonThread_1_io_output_payload_stateSize;
  wire       [7:0]    poseidonThread_1_io_output_payload_stateID;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_0;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_1;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_2;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_3;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_4;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_5;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_6;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_7;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_8;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_9;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_10;
  wire       [254:0]  poseidonThread_1_io_output_payload_stateElements_11;
  wire                demuxInst_io_input_ready;
  wire                demuxInst_io_output0_valid;
  wire                demuxInst_io_output0_payload_isFull;
  wire       [2:0]    demuxInst_io_output0_payload_fullRound;
  wire       [5:0]    demuxInst_io_output0_payload_partialRound;
  wire       [3:0]    demuxInst_io_output0_payload_stateSize;
  wire       [7:0]    demuxInst_io_output0_payload_stateID;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_0;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_1;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_2;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_3;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_4;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_5;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_6;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_7;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_8;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_9;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_10;
  wire       [254:0]  demuxInst_io_output0_payload_stateElements_11;
  wire                demuxInst_io_output1_valid;
  wire       [7:0]    demuxInst_io_output1_payload_stateID;
  wire       [254:0]  demuxInst_io_output1_payload_stateElement;
  wire                bundleFifo_1_io_push_ready;
  wire                bundleFifo_1_io_pop_valid;
  wire                bundleFifo_1_io_pop_payload_isFull;
  wire       [2:0]    bundleFifo_1_io_pop_payload_fullRound;
  wire       [5:0]    bundleFifo_1_io_pop_payload_partialRound;
  wire       [3:0]    bundleFifo_1_io_pop_payload_stateSize;
  wire       [7:0]    bundleFifo_1_io_pop_payload_stateID;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_0;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_1;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_2;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_3;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_4;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_5;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_6;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_7;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_8;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_9;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_10;
  wire       [254:0]  bundleFifo_1_io_pop_payload_stateElements_11;
  wire                loopbackBuffer_valid;
  wire                loopbackBuffer_ready;
  wire                loopbackBuffer_payload_isFull;
  wire       [2:0]    loopbackBuffer_payload_fullRound;
  wire       [5:0]    loopbackBuffer_payload_partialRound;
  wire       [3:0]    loopbackBuffer_payload_stateSize;
  wire       [7:0]    loopbackBuffer_payload_stateID;
  wire       [254:0]  loopbackBuffer_payload_stateElements_0;
  wire       [254:0]  loopbackBuffer_payload_stateElements_1;
  wire       [254:0]  loopbackBuffer_payload_stateElements_2;
  wire       [254:0]  loopbackBuffer_payload_stateElements_3;
  wire       [254:0]  loopbackBuffer_payload_stateElements_4;
  wire       [254:0]  loopbackBuffer_payload_stateElements_5;
  wire       [254:0]  loopbackBuffer_payload_stateElements_6;
  wire       [254:0]  loopbackBuffer_payload_stateElements_7;
  wire       [254:0]  loopbackBuffer_payload_stateElements_8;
  wire       [254:0]  loopbackBuffer_payload_stateElements_9;
  wire       [254:0]  loopbackBuffer_payload_stateElements_10;
  wire       [254:0]  loopbackBuffer_payload_stateElements_11;
  wire                preRoundConstStage_input_valid;
  wire                preRoundConstStage_input_payload_isFull;
  wire       [2:0]    preRoundConstStage_input_payload_fullRound;
  wire       [5:0]    preRoundConstStage_input_payload_partialRound;
  wire       [3:0]    preRoundConstStage_input_payload_stateIndex;
  wire       [3:0]    preRoundConstStage_input_payload_stateSize;
  wire       [7:0]    preRoundConstStage_input_payload_stateID;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_0;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_1;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_2;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_3;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_4;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_5;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_6;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_7;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_8;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_9;
  wire       [254:0]  preRoundConstStage_input_payload_stateElements_10;
  wire       [254:0]  preRoundConstStage_input_payload_stateElement;
  wire                preRoundConstStage_adderInput_valid;
  wire       [254:0]  preRoundConstStage_adderInput_payload_op1;
  wire       [254:0]  preRoundConstStage_adderInput_payload_op2;
  reg                 preRoundConstStage_input_payload_delay_1_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_1_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_1_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_1_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_1_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_1_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_1_stateElement;
  reg                 preRoundConstStage_input_payload_delay_2_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_2_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_2_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_2_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_2_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_2_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_2_stateElement;
  reg                 preRoundConstStage_input_payload_delay_3_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_3_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_3_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_3_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_3_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_3_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_3_stateElement;
  reg                 preRoundConstStage_input_payload_delay_4_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_4_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_4_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_4_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_4_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_4_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_4_stateElement;
  reg                 preRoundConstStage_input_payload_delay_5_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_5_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_5_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_5_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_5_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_5_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_5_stateElement;
  reg                 preRoundConstStage_input_payload_delay_6_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_6_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_6_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_6_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_6_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_6_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_6_stateElement;
  reg                 preRoundConstStage_input_payload_delay_7_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_7_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_7_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_7_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_7_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_7_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_7_stateElement;
  reg                 preRoundConstStage_input_payload_delay_8_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_8_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_8_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_8_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_8_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_8_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_8_stateElement;
  reg                 preRoundConstStage_input_payload_delay_9_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_9_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_9_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_9_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_9_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_9_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_9_stateElement;
  reg                 preRoundConstStage_input_payload_delay_10_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_10_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_10_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_10_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_10_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_10_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_10_stateElement;
  reg                 preRoundConstStage_input_payload_delay_11_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_11_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_11_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_11_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_11_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_11_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_11_stateElement;
  reg                 preRoundConstStage_input_payload_delay_12_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_12_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_12_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_12_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_12_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_12_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_12_stateElement;
  reg                 preRoundConstStage_input_payload_delay_13_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_13_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_13_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_13_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_13_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_13_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_13_stateElement;
  reg                 preRoundConstStage_input_payload_delay_14_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_14_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_14_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_14_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_14_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_14_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_14_stateElement;
  reg                 preRoundConstStage_input_payload_delay_15_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_15_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_15_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_15_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_15_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_15_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_15_stateElement;
  reg                 preRoundConstStage_input_payload_delay_16_isFull;
  reg        [2:0]    preRoundConstStage_input_payload_delay_16_fullRound;
  reg        [5:0]    preRoundConstStage_input_payload_delay_16_partialRound;
  reg        [3:0]    preRoundConstStage_input_payload_delay_16_stateIndex;
  reg        [3:0]    preRoundConstStage_input_payload_delay_16_stateSize;
  reg        [7:0]    preRoundConstStage_input_payload_delay_16_stateID;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_0;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_1;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_2;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_3;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_4;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_5;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_6;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_7;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_8;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_9;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElements_10;
  reg        [254:0]  preRoundConstStage_input_payload_delay_16_stateElement;
  reg                 preRoundConstStage_addContextDelayed_isFull;
  reg        [2:0]    preRoundConstStage_addContextDelayed_fullRound;
  reg        [5:0]    preRoundConstStage_addContextDelayed_partialRound;
  reg        [3:0]    preRoundConstStage_addContextDelayed_stateIndex;
  reg        [3:0]    preRoundConstStage_addContextDelayed_stateSize;
  reg        [7:0]    preRoundConstStage_addContextDelayed_stateID;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_0;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_1;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_2;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_3;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_4;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_5;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_6;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_7;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_8;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_9;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElements_10;
  reg        [254:0]  preRoundConstStage_addContextDelayed_stateElement;
  wire                preRoundConstStage_output_valid;
  wire                preRoundConstStage_output_payload_isFull;
  wire       [2:0]    preRoundConstStage_output_payload_fullRound;
  wire       [5:0]    preRoundConstStage_output_payload_partialRound;
  wire       [3:0]    preRoundConstStage_output_payload_stateIndex;
  wire       [3:0]    preRoundConstStage_output_payload_stateSize;
  wire       [7:0]    preRoundConstStage_output_payload_stateID;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_0;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_1;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_2;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_3;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_4;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_5;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_6;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_7;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_8;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_9;
  wire       [254:0]  preRoundConstStage_output_payload_stateElements_10;
  reg        [254:0]  preRoundConstStage_output_payload_stateElement;
  wire                when_PoseidonTopLevel_l173;
  wire                poseidonThread_1_io_output_toStream_valid;
  wire                poseidonThread_1_io_output_toStream_ready;
  wire                poseidonThread_1_io_output_toStream_payload_isFull;
  wire       [2:0]    poseidonThread_1_io_output_toStream_payload_fullRound;
  wire       [5:0]    poseidonThread_1_io_output_toStream_payload_partialRound;
  wire       [3:0]    poseidonThread_1_io_output_toStream_payload_stateSize;
  wire       [7:0]    poseidonThread_1_io_output_toStream_payload_stateID;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_0;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_1;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_2;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_3;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_4;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_5;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_6;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_7;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_8;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_9;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_10;
  wire       [254:0]  poseidonThread_1_io_output_toStream_payload_stateElements_11;
  wire                demuxInst_io_output0_s2mPipe_valid;
  reg                 demuxInst_io_output0_s2mPipe_ready;
  wire                demuxInst_io_output0_s2mPipe_payload_isFull;
  wire       [2:0]    demuxInst_io_output0_s2mPipe_payload_fullRound;
  wire       [5:0]    demuxInst_io_output0_s2mPipe_payload_partialRound;
  wire       [3:0]    demuxInst_io_output0_s2mPipe_payload_stateSize;
  wire       [7:0]    demuxInst_io_output0_s2mPipe_payload_stateID;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_0;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_1;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_2;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_3;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_4;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_5;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_6;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_7;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_8;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_9;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_10;
  wire       [254:0]  demuxInst_io_output0_s2mPipe_payload_stateElements_11;
  reg                 demuxInst_io_output0_rValid;
  reg                 demuxInst_io_output0_rData_isFull;
  reg        [2:0]    demuxInst_io_output0_rData_fullRound;
  reg        [5:0]    demuxInst_io_output0_rData_partialRound;
  reg        [3:0]    demuxInst_io_output0_rData_stateSize;
  reg        [7:0]    demuxInst_io_output0_rData_stateID;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_0;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_1;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_2;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_3;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_4;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_5;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_6;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_7;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_8;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_9;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_10;
  reg        [254:0]  demuxInst_io_output0_rData_stateElements_11;
  wire                loopback_valid;
  wire                loopback_ready;
  wire                loopback_payload_isFull;
  wire       [2:0]    loopback_payload_fullRound;
  wire       [5:0]    loopback_payload_partialRound;
  wire       [3:0]    loopback_payload_stateSize;
  wire       [7:0]    loopback_payload_stateID;
  wire       [254:0]  loopback_payload_stateElements_0;
  wire       [254:0]  loopback_payload_stateElements_1;
  wire       [254:0]  loopback_payload_stateElements_2;
  wire       [254:0]  loopback_payload_stateElements_3;
  wire       [254:0]  loopback_payload_stateElements_4;
  wire       [254:0]  loopback_payload_stateElements_5;
  wire       [254:0]  loopback_payload_stateElements_6;
  wire       [254:0]  loopback_payload_stateElements_7;
  wire       [254:0]  loopback_payload_stateElements_8;
  wire       [254:0]  loopback_payload_stateElements_9;
  wire       [254:0]  loopback_payload_stateElements_10;
  wire       [254:0]  loopback_payload_stateElements_11;
  reg                 demuxInst_io_output0_s2mPipe_rValid;
  reg                 demuxInst_io_output0_s2mPipe_rData_isFull;
  reg        [2:0]    demuxInst_io_output0_s2mPipe_rData_fullRound;
  reg        [5:0]    demuxInst_io_output0_s2mPipe_rData_partialRound;
  reg        [3:0]    demuxInst_io_output0_s2mPipe_rData_stateSize;
  reg        [7:0]    demuxInst_io_output0_s2mPipe_rData_stateID;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_0;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_1;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_2;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_3;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_4;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_5;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_6;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_7;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_8;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_9;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_10;
  reg        [254:0]  demuxInst_io_output0_s2mPipe_rData_stateElements_11;
  wire                when_Stream_l342;
  wire                demuxInst_io_output1_m2sPipe_valid;
  wire                demuxInst_io_output1_m2sPipe_ready;
  wire       [7:0]    demuxInst_io_output1_m2sPipe_payload_stateID;
  wire       [254:0]  demuxInst_io_output1_m2sPipe_payload_stateElement;
  reg                 demuxInst_io_output1_rValid;
  reg        [7:0]    demuxInst_io_output1_rData_stateID;
  reg        [254:0]  demuxInst_io_output1_rData_stateElement;
  wire                when_Stream_l342_1;

  StreamArbiter streamArbiter_2 (
    .io_inputs_0_valid                       (loopbackBuffer_valid                                       ), //i
    .io_inputs_0_ready                       (streamArbiter_2_io_inputs_0_ready                          ), //o
    .io_inputs_0_payload_isFull              (loopbackBuffer_payload_isFull                              ), //i
    .io_inputs_0_payload_fullRound           (loopbackBuffer_payload_fullRound[2:0]                      ), //i
    .io_inputs_0_payload_partialRound        (loopbackBuffer_payload_partialRound[5:0]                   ), //i
    .io_inputs_0_payload_stateSize           (loopbackBuffer_payload_stateSize[3:0]                      ), //i
    .io_inputs_0_payload_stateID             (loopbackBuffer_payload_stateID[7:0]                        ), //i
    .io_inputs_0_payload_stateElements_0     (loopbackBuffer_payload_stateElements_0[254:0]              ), //i
    .io_inputs_0_payload_stateElements_1     (loopbackBuffer_payload_stateElements_1[254:0]              ), //i
    .io_inputs_0_payload_stateElements_2     (loopbackBuffer_payload_stateElements_2[254:0]              ), //i
    .io_inputs_0_payload_stateElements_3     (loopbackBuffer_payload_stateElements_3[254:0]              ), //i
    .io_inputs_0_payload_stateElements_4     (loopbackBuffer_payload_stateElements_4[254:0]              ), //i
    .io_inputs_0_payload_stateElements_5     (loopbackBuffer_payload_stateElements_5[254:0]              ), //i
    .io_inputs_0_payload_stateElements_6     (loopbackBuffer_payload_stateElements_6[254:0]              ), //i
    .io_inputs_0_payload_stateElements_7     (loopbackBuffer_payload_stateElements_7[254:0]              ), //i
    .io_inputs_0_payload_stateElements_8     (loopbackBuffer_payload_stateElements_8[254:0]              ), //i
    .io_inputs_0_payload_stateElements_9     (loopbackBuffer_payload_stateElements_9[254:0]              ), //i
    .io_inputs_0_payload_stateElements_10    (loopbackBuffer_payload_stateElements_10[254:0]             ), //i
    .io_inputs_0_payload_stateElements_11    (loopbackBuffer_payload_stateElements_11[254:0]             ), //i
    .io_inputs_1_valid                       (io_input_valid                                             ), //i
    .io_inputs_1_ready                       (streamArbiter_2_io_inputs_1_ready                          ), //o
    .io_inputs_1_payload_isFull              (io_input_payload_isFull                                    ), //i
    .io_inputs_1_payload_fullRound           (io_input_payload_fullRound[2:0]                            ), //i
    .io_inputs_1_payload_partialRound        (io_input_payload_partialRound[5:0]                         ), //i
    .io_inputs_1_payload_stateSize           (io_input_payload_stateSize[3:0]                            ), //i
    .io_inputs_1_payload_stateID             (io_input_payload_stateID[7:0]                              ), //i
    .io_inputs_1_payload_stateElements_0     (io_input_payload_stateElements_0[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_1     (io_input_payload_stateElements_1[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_2     (io_input_payload_stateElements_2[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_3     (io_input_payload_stateElements_3[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_4     (io_input_payload_stateElements_4[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_5     (io_input_payload_stateElements_5[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_6     (io_input_payload_stateElements_6[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_7     (io_input_payload_stateElements_7[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_8     (io_input_payload_stateElements_8[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_9     (io_input_payload_stateElements_9[254:0]                    ), //i
    .io_inputs_1_payload_stateElements_10    (io_input_payload_stateElements_10[254:0]                   ), //i
    .io_inputs_1_payload_stateElements_11    (io_input_payload_stateElements_11[254:0]                   ), //i
    .io_output_valid                         (streamArbiter_2_io_output_valid                            ), //o
    .io_output_ready                         (poseidonSerializer_1_io_input_ready                        ), //i
    .io_output_payload_isFull                (streamArbiter_2_io_output_payload_isFull                   ), //o
    .io_output_payload_fullRound             (streamArbiter_2_io_output_payload_fullRound[2:0]           ), //o
    .io_output_payload_partialRound          (streamArbiter_2_io_output_payload_partialRound[5:0]        ), //o
    .io_output_payload_stateSize             (streamArbiter_2_io_output_payload_stateSize[3:0]           ), //o
    .io_output_payload_stateID               (streamArbiter_2_io_output_payload_stateID[7:0]             ), //o
    .io_output_payload_stateElements_0       (streamArbiter_2_io_output_payload_stateElements_0[254:0]   ), //o
    .io_output_payload_stateElements_1       (streamArbiter_2_io_output_payload_stateElements_1[254:0]   ), //o
    .io_output_payload_stateElements_2       (streamArbiter_2_io_output_payload_stateElements_2[254:0]   ), //o
    .io_output_payload_stateElements_3       (streamArbiter_2_io_output_payload_stateElements_3[254:0]   ), //o
    .io_output_payload_stateElements_4       (streamArbiter_2_io_output_payload_stateElements_4[254:0]   ), //o
    .io_output_payload_stateElements_5       (streamArbiter_2_io_output_payload_stateElements_5[254:0]   ), //o
    .io_output_payload_stateElements_6       (streamArbiter_2_io_output_payload_stateElements_6[254:0]   ), //o
    .io_output_payload_stateElements_7       (streamArbiter_2_io_output_payload_stateElements_7[254:0]   ), //o
    .io_output_payload_stateElements_8       (streamArbiter_2_io_output_payload_stateElements_8[254:0]   ), //o
    .io_output_payload_stateElements_9       (streamArbiter_2_io_output_payload_stateElements_9[254:0]   ), //o
    .io_output_payload_stateElements_10      (streamArbiter_2_io_output_payload_stateElements_10[254:0]  ), //o
    .io_output_payload_stateElements_11      (streamArbiter_2_io_output_payload_stateElements_11[254:0]  ), //o
    .io_chosen                               (streamArbiter_2_io_chosen                                  ), //o
    .io_chosenOH                             (streamArbiter_2_io_chosenOH[1:0]                           ), //o
    .clk                                     (clk                                                        ), //i
    .resetn                                  (resetn                                                     )  //i
  );
  PoseidonSerializer poseidonSerializer_1 (
    .io_input_valid                        (streamArbiter_2_io_output_valid                                 ), //i
    .io_input_ready                        (poseidonSerializer_1_io_input_ready                             ), //o
    .io_input_payload_isFull               (streamArbiter_2_io_output_payload_isFull                        ), //i
    .io_input_payload_fullRound            (streamArbiter_2_io_output_payload_fullRound[2:0]                ), //i
    .io_input_payload_partialRound         (streamArbiter_2_io_output_payload_partialRound[5:0]             ), //i
    .io_input_payload_stateSize            (streamArbiter_2_io_output_payload_stateSize[3:0]                ), //i
    .io_input_payload_stateID              (streamArbiter_2_io_output_payload_stateID[7:0]                  ), //i
    .io_input_payload_stateElements_0      (streamArbiter_2_io_output_payload_stateElements_0[254:0]        ), //i
    .io_input_payload_stateElements_1      (streamArbiter_2_io_output_payload_stateElements_1[254:0]        ), //i
    .io_input_payload_stateElements_2      (streamArbiter_2_io_output_payload_stateElements_2[254:0]        ), //i
    .io_input_payload_stateElements_3      (streamArbiter_2_io_output_payload_stateElements_3[254:0]        ), //i
    .io_input_payload_stateElements_4      (streamArbiter_2_io_output_payload_stateElements_4[254:0]        ), //i
    .io_input_payload_stateElements_5      (streamArbiter_2_io_output_payload_stateElements_5[254:0]        ), //i
    .io_input_payload_stateElements_6      (streamArbiter_2_io_output_payload_stateElements_6[254:0]        ), //i
    .io_input_payload_stateElements_7      (streamArbiter_2_io_output_payload_stateElements_7[254:0]        ), //i
    .io_input_payload_stateElements_8      (streamArbiter_2_io_output_payload_stateElements_8[254:0]        ), //i
    .io_input_payload_stateElements_9      (streamArbiter_2_io_output_payload_stateElements_9[254:0]        ), //i
    .io_input_payload_stateElements_10     (streamArbiter_2_io_output_payload_stateElements_10[254:0]       ), //i
    .io_input_payload_stateElements_11     (streamArbiter_2_io_output_payload_stateElements_11[254:0]       ), //i
    .io_output_valid                       (poseidonSerializer_1_io_output_valid                            ), //o
    .io_output_ready                       (1'b1                                                            ), //i
    .io_output_payload_isFull              (poseidonSerializer_1_io_output_payload_isFull                   ), //o
    .io_output_payload_fullRound           (poseidonSerializer_1_io_output_payload_fullRound[2:0]           ), //o
    .io_output_payload_partialRound        (poseidonSerializer_1_io_output_payload_partialRound[5:0]        ), //o
    .io_output_payload_stateIndex          (poseidonSerializer_1_io_output_payload_stateIndex[3:0]          ), //o
    .io_output_payload_stateSize           (poseidonSerializer_1_io_output_payload_stateSize[3:0]           ), //o
    .io_output_payload_stateID             (poseidonSerializer_1_io_output_payload_stateID[7:0]             ), //o
    .io_output_payload_stateElements_0     (poseidonSerializer_1_io_output_payload_stateElements_0[254:0]   ), //o
    .io_output_payload_stateElements_1     (poseidonSerializer_1_io_output_payload_stateElements_1[254:0]   ), //o
    .io_output_payload_stateElements_2     (poseidonSerializer_1_io_output_payload_stateElements_2[254:0]   ), //o
    .io_output_payload_stateElements_3     (poseidonSerializer_1_io_output_payload_stateElements_3[254:0]   ), //o
    .io_output_payload_stateElements_4     (poseidonSerializer_1_io_output_payload_stateElements_4[254:0]   ), //o
    .io_output_payload_stateElements_5     (poseidonSerializer_1_io_output_payload_stateElements_5[254:0]   ), //o
    .io_output_payload_stateElements_6     (poseidonSerializer_1_io_output_payload_stateElements_6[254:0]   ), //o
    .io_output_payload_stateElements_7     (poseidonSerializer_1_io_output_payload_stateElements_7[254:0]   ), //o
    .io_output_payload_stateElements_8     (poseidonSerializer_1_io_output_payload_stateElements_8[254:0]   ), //o
    .io_output_payload_stateElements_9     (poseidonSerializer_1_io_output_payload_stateElements_9[254:0]   ), //o
    .io_output_payload_stateElements_10    (poseidonSerializer_1_io_output_payload_stateElements_10[254:0]  ), //o
    .io_output_payload_stateElement        (poseidonSerializer_1_io_output_payload_stateElement[254:0]      ), //o
    .clk                                   (clk                                                             ), //i
    .resetn                                (resetn                                                          )  //i
  );
  PreRoundConstantMem preRoundConstantMem_1 (
    .io_stateSize      (preRoundConstStage_input_payload_stateSize[3:0]   ), //i
    .io_stateIndex     (preRoundConstStage_input_payload_stateIndex[3:0]  ), //i
    .io_preConstant    (preRoundConstantMem_1_io_preConstant[254:0]       )  //o
  );
  ModularAdderFlow_1 preRoundConstStage_adderInst (
    .io_input_valid           (preRoundConstStage_adderInput_valid                        ), //i
    .io_input_payload_op1     (preRoundConstStage_adderInput_payload_op1[254:0]           ), //i
    .io_input_payload_op2     (preRoundConstStage_adderInput_payload_op2[254:0]           ), //i
    .io_output_valid          (preRoundConstStage_adderInst_io_output_valid               ), //o
    .io_output_payload_res    (preRoundConstStage_adderInst_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                        ), //i
    .resetn                   (resetn                                                     )  //i
  );
  PoseidonThread poseidonThread_1 (
    .io_input_valid                        (preRoundConstStage_output_valid                             ), //i
    .io_input_payload_isFull               (preRoundConstStage_output_payload_isFull                    ), //i
    .io_input_payload_fullRound            (preRoundConstStage_output_payload_fullRound[2:0]            ), //i
    .io_input_payload_partialRound         (preRoundConstStage_output_payload_partialRound[5:0]         ), //i
    .io_input_payload_stateIndex           (preRoundConstStage_output_payload_stateIndex[3:0]           ), //i
    .io_input_payload_stateSize            (preRoundConstStage_output_payload_stateSize[3:0]            ), //i
    .io_input_payload_stateID              (preRoundConstStage_output_payload_stateID[7:0]              ), //i
    .io_input_payload_stateElements_0      (preRoundConstStage_output_payload_stateElements_0[254:0]    ), //i
    .io_input_payload_stateElements_1      (preRoundConstStage_output_payload_stateElements_1[254:0]    ), //i
    .io_input_payload_stateElements_2      (preRoundConstStage_output_payload_stateElements_2[254:0]    ), //i
    .io_input_payload_stateElements_3      (preRoundConstStage_output_payload_stateElements_3[254:0]    ), //i
    .io_input_payload_stateElements_4      (preRoundConstStage_output_payload_stateElements_4[254:0]    ), //i
    .io_input_payload_stateElements_5      (preRoundConstStage_output_payload_stateElements_5[254:0]    ), //i
    .io_input_payload_stateElements_6      (preRoundConstStage_output_payload_stateElements_6[254:0]    ), //i
    .io_input_payload_stateElements_7      (preRoundConstStage_output_payload_stateElements_7[254:0]    ), //i
    .io_input_payload_stateElements_8      (preRoundConstStage_output_payload_stateElements_8[254:0]    ), //i
    .io_input_payload_stateElements_9      (preRoundConstStage_output_payload_stateElements_9[254:0]    ), //i
    .io_input_payload_stateElements_10     (preRoundConstStage_output_payload_stateElements_10[254:0]   ), //i
    .io_input_payload_stateElement         (preRoundConstStage_output_payload_stateElement[254:0]       ), //i
    .io_output_valid                       (poseidonThread_1_io_output_valid                            ), //o
    .io_output_payload_isFull              (poseidonThread_1_io_output_payload_isFull                   ), //o
    .io_output_payload_fullRound           (poseidonThread_1_io_output_payload_fullRound[2:0]           ), //o
    .io_output_payload_partialRound        (poseidonThread_1_io_output_payload_partialRound[5:0]        ), //o
    .io_output_payload_stateSize           (poseidonThread_1_io_output_payload_stateSize[3:0]           ), //o
    .io_output_payload_stateID             (poseidonThread_1_io_output_payload_stateID[7:0]             ), //o
    .io_output_payload_stateElements_0     (poseidonThread_1_io_output_payload_stateElements_0[254:0]   ), //o
    .io_output_payload_stateElements_1     (poseidonThread_1_io_output_payload_stateElements_1[254:0]   ), //o
    .io_output_payload_stateElements_2     (poseidonThread_1_io_output_payload_stateElements_2[254:0]   ), //o
    .io_output_payload_stateElements_3     (poseidonThread_1_io_output_payload_stateElements_3[254:0]   ), //o
    .io_output_payload_stateElements_4     (poseidonThread_1_io_output_payload_stateElements_4[254:0]   ), //o
    .io_output_payload_stateElements_5     (poseidonThread_1_io_output_payload_stateElements_5[254:0]   ), //o
    .io_output_payload_stateElements_6     (poseidonThread_1_io_output_payload_stateElements_6[254:0]   ), //o
    .io_output_payload_stateElements_7     (poseidonThread_1_io_output_payload_stateElements_7[254:0]   ), //o
    .io_output_payload_stateElements_8     (poseidonThread_1_io_output_payload_stateElements_8[254:0]   ), //o
    .io_output_payload_stateElements_9     (poseidonThread_1_io_output_payload_stateElements_9[254:0]   ), //o
    .io_output_payload_stateElements_10    (poseidonThread_1_io_output_payload_stateElements_10[254:0]  ), //o
    .io_output_payload_stateElements_11    (poseidonThread_1_io_output_payload_stateElements_11[254:0]  ), //o
    .clk                                   (clk                                                         ), //i
    .resetn                                (resetn                                                      )  //i
  );
  LoopbackDeMux demuxInst (
    .io_input_valid                         (poseidonThread_1_io_output_toStream_valid                            ), //i
    .io_input_ready                         (demuxInst_io_input_ready                                             ), //o
    .io_input_payload_isFull                (poseidonThread_1_io_output_toStream_payload_isFull                   ), //i
    .io_input_payload_fullRound             (poseidonThread_1_io_output_toStream_payload_fullRound[2:0]           ), //i
    .io_input_payload_partialRound          (poseidonThread_1_io_output_toStream_payload_partialRound[5:0]        ), //i
    .io_input_payload_stateSize             (poseidonThread_1_io_output_toStream_payload_stateSize[3:0]           ), //i
    .io_input_payload_stateID               (poseidonThread_1_io_output_toStream_payload_stateID[7:0]             ), //i
    .io_input_payload_stateElements_0       (poseidonThread_1_io_output_toStream_payload_stateElements_0[254:0]   ), //i
    .io_input_payload_stateElements_1       (poseidonThread_1_io_output_toStream_payload_stateElements_1[254:0]   ), //i
    .io_input_payload_stateElements_2       (poseidonThread_1_io_output_toStream_payload_stateElements_2[254:0]   ), //i
    .io_input_payload_stateElements_3       (poseidonThread_1_io_output_toStream_payload_stateElements_3[254:0]   ), //i
    .io_input_payload_stateElements_4       (poseidonThread_1_io_output_toStream_payload_stateElements_4[254:0]   ), //i
    .io_input_payload_stateElements_5       (poseidonThread_1_io_output_toStream_payload_stateElements_5[254:0]   ), //i
    .io_input_payload_stateElements_6       (poseidonThread_1_io_output_toStream_payload_stateElements_6[254:0]   ), //i
    .io_input_payload_stateElements_7       (poseidonThread_1_io_output_toStream_payload_stateElements_7[254:0]   ), //i
    .io_input_payload_stateElements_8       (poseidonThread_1_io_output_toStream_payload_stateElements_8[254:0]   ), //i
    .io_input_payload_stateElements_9       (poseidonThread_1_io_output_toStream_payload_stateElements_9[254:0]   ), //i
    .io_input_payload_stateElements_10      (poseidonThread_1_io_output_toStream_payload_stateElements_10[254:0]  ), //i
    .io_input_payload_stateElements_11      (poseidonThread_1_io_output_toStream_payload_stateElements_11[254:0]  ), //i
    .io_output0_valid                       (demuxInst_io_output0_valid                                           ), //o
    .io_output0_ready                       (demuxInst_io_output0_ready                                           ), //i
    .io_output0_payload_isFull              (demuxInst_io_output0_payload_isFull                                  ), //o
    .io_output0_payload_fullRound           (demuxInst_io_output0_payload_fullRound[2:0]                          ), //o
    .io_output0_payload_partialRound        (demuxInst_io_output0_payload_partialRound[5:0]                       ), //o
    .io_output0_payload_stateSize           (demuxInst_io_output0_payload_stateSize[3:0]                          ), //o
    .io_output0_payload_stateID             (demuxInst_io_output0_payload_stateID[7:0]                            ), //o
    .io_output0_payload_stateElements_0     (demuxInst_io_output0_payload_stateElements_0[254:0]                  ), //o
    .io_output0_payload_stateElements_1     (demuxInst_io_output0_payload_stateElements_1[254:0]                  ), //o
    .io_output0_payload_stateElements_2     (demuxInst_io_output0_payload_stateElements_2[254:0]                  ), //o
    .io_output0_payload_stateElements_3     (demuxInst_io_output0_payload_stateElements_3[254:0]                  ), //o
    .io_output0_payload_stateElements_4     (demuxInst_io_output0_payload_stateElements_4[254:0]                  ), //o
    .io_output0_payload_stateElements_5     (demuxInst_io_output0_payload_stateElements_5[254:0]                  ), //o
    .io_output0_payload_stateElements_6     (demuxInst_io_output0_payload_stateElements_6[254:0]                  ), //o
    .io_output0_payload_stateElements_7     (demuxInst_io_output0_payload_stateElements_7[254:0]                  ), //o
    .io_output0_payload_stateElements_8     (demuxInst_io_output0_payload_stateElements_8[254:0]                  ), //o
    .io_output0_payload_stateElements_9     (demuxInst_io_output0_payload_stateElements_9[254:0]                  ), //o
    .io_output0_payload_stateElements_10    (demuxInst_io_output0_payload_stateElements_10[254:0]                 ), //o
    .io_output0_payload_stateElements_11    (demuxInst_io_output0_payload_stateElements_11[254:0]                 ), //o
    .io_output1_valid                       (demuxInst_io_output1_valid                                           ), //o
    .io_output1_ready                       (demuxInst_io_output1_ready                                           ), //i
    .io_output1_payload_stateID             (demuxInst_io_output1_payload_stateID[7:0]                            ), //o
    .io_output1_payload_stateElement        (demuxInst_io_output1_payload_stateElement[254:0]                     )  //o
  );
  BundleFifo bundleFifo_1 (
    .io_push_valid                       (loopback_valid                                       ), //i
    .io_push_ready                       (bundleFifo_1_io_push_ready                           ), //o
    .io_push_payload_isFull              (loopback_payload_isFull                              ), //i
    .io_push_payload_fullRound           (loopback_payload_fullRound[2:0]                      ), //i
    .io_push_payload_partialRound        (loopback_payload_partialRound[5:0]                   ), //i
    .io_push_payload_stateSize           (loopback_payload_stateSize[3:0]                      ), //i
    .io_push_payload_stateID             (loopback_payload_stateID[7:0]                        ), //i
    .io_push_payload_stateElements_0     (loopback_payload_stateElements_0[254:0]              ), //i
    .io_push_payload_stateElements_1     (loopback_payload_stateElements_1[254:0]              ), //i
    .io_push_payload_stateElements_2     (loopback_payload_stateElements_2[254:0]              ), //i
    .io_push_payload_stateElements_3     (loopback_payload_stateElements_3[254:0]              ), //i
    .io_push_payload_stateElements_4     (loopback_payload_stateElements_4[254:0]              ), //i
    .io_push_payload_stateElements_5     (loopback_payload_stateElements_5[254:0]              ), //i
    .io_push_payload_stateElements_6     (loopback_payload_stateElements_6[254:0]              ), //i
    .io_push_payload_stateElements_7     (loopback_payload_stateElements_7[254:0]              ), //i
    .io_push_payload_stateElements_8     (loopback_payload_stateElements_8[254:0]              ), //i
    .io_push_payload_stateElements_9     (loopback_payload_stateElements_9[254:0]              ), //i
    .io_push_payload_stateElements_10    (loopback_payload_stateElements_10[254:0]             ), //i
    .io_push_payload_stateElements_11    (loopback_payload_stateElements_11[254:0]             ), //i
    .io_pop_valid                        (bundleFifo_1_io_pop_valid                            ), //o
    .io_pop_ready                        (loopbackBuffer_ready                                 ), //i
    .io_pop_payload_isFull               (bundleFifo_1_io_pop_payload_isFull                   ), //o
    .io_pop_payload_fullRound            (bundleFifo_1_io_pop_payload_fullRound[2:0]           ), //o
    .io_pop_payload_partialRound         (bundleFifo_1_io_pop_payload_partialRound[5:0]        ), //o
    .io_pop_payload_stateSize            (bundleFifo_1_io_pop_payload_stateSize[3:0]           ), //o
    .io_pop_payload_stateID              (bundleFifo_1_io_pop_payload_stateID[7:0]             ), //o
    .io_pop_payload_stateElements_0      (bundleFifo_1_io_pop_payload_stateElements_0[254:0]   ), //o
    .io_pop_payload_stateElements_1      (bundleFifo_1_io_pop_payload_stateElements_1[254:0]   ), //o
    .io_pop_payload_stateElements_2      (bundleFifo_1_io_pop_payload_stateElements_2[254:0]   ), //o
    .io_pop_payload_stateElements_3      (bundleFifo_1_io_pop_payload_stateElements_3[254:0]   ), //o
    .io_pop_payload_stateElements_4      (bundleFifo_1_io_pop_payload_stateElements_4[254:0]   ), //o
    .io_pop_payload_stateElements_5      (bundleFifo_1_io_pop_payload_stateElements_5[254:0]   ), //o
    .io_pop_payload_stateElements_6      (bundleFifo_1_io_pop_payload_stateElements_6[254:0]   ), //o
    .io_pop_payload_stateElements_7      (bundleFifo_1_io_pop_payload_stateElements_7[254:0]   ), //o
    .io_pop_payload_stateElements_8      (bundleFifo_1_io_pop_payload_stateElements_8[254:0]   ), //o
    .io_pop_payload_stateElements_9      (bundleFifo_1_io_pop_payload_stateElements_9[254:0]   ), //o
    .io_pop_payload_stateElements_10     (bundleFifo_1_io_pop_payload_stateElements_10[254:0]  ), //o
    .io_pop_payload_stateElements_11     (bundleFifo_1_io_pop_payload_stateElements_11[254:0]  ), //o
    .clk                                 (clk                                                  ), //i
    .resetn                              (resetn                                               )  //i
  );
  assign loopbackBuffer_ready = streamArbiter_2_io_inputs_0_ready;
  assign io_input_ready = streamArbiter_2_io_inputs_1_ready;
  assign preRoundConstStage_input_valid = poseidonSerializer_1_io_output_valid;
  assign preRoundConstStage_input_payload_isFull = poseidonSerializer_1_io_output_payload_isFull;
  assign preRoundConstStage_input_payload_fullRound = poseidonSerializer_1_io_output_payload_fullRound;
  assign preRoundConstStage_input_payload_partialRound = poseidonSerializer_1_io_output_payload_partialRound;
  assign preRoundConstStage_input_payload_stateIndex = poseidonSerializer_1_io_output_payload_stateIndex;
  assign preRoundConstStage_input_payload_stateSize = poseidonSerializer_1_io_output_payload_stateSize;
  assign preRoundConstStage_input_payload_stateID = poseidonSerializer_1_io_output_payload_stateID;
  assign preRoundConstStage_input_payload_stateElements_0 = poseidonSerializer_1_io_output_payload_stateElements_0;
  assign preRoundConstStage_input_payload_stateElements_1 = poseidonSerializer_1_io_output_payload_stateElements_1;
  assign preRoundConstStage_input_payload_stateElements_2 = poseidonSerializer_1_io_output_payload_stateElements_2;
  assign preRoundConstStage_input_payload_stateElements_3 = poseidonSerializer_1_io_output_payload_stateElements_3;
  assign preRoundConstStage_input_payload_stateElements_4 = poseidonSerializer_1_io_output_payload_stateElements_4;
  assign preRoundConstStage_input_payload_stateElements_5 = poseidonSerializer_1_io_output_payload_stateElements_5;
  assign preRoundConstStage_input_payload_stateElements_6 = poseidonSerializer_1_io_output_payload_stateElements_6;
  assign preRoundConstStage_input_payload_stateElements_7 = poseidonSerializer_1_io_output_payload_stateElements_7;
  assign preRoundConstStage_input_payload_stateElements_8 = poseidonSerializer_1_io_output_payload_stateElements_8;
  assign preRoundConstStage_input_payload_stateElements_9 = poseidonSerializer_1_io_output_payload_stateElements_9;
  assign preRoundConstStage_input_payload_stateElements_10 = poseidonSerializer_1_io_output_payload_stateElements_10;
  assign preRoundConstStage_input_payload_stateElement = poseidonSerializer_1_io_output_payload_stateElement;
  assign preRoundConstStage_adderInput_valid = preRoundConstStage_input_valid;
  assign preRoundConstStage_adderInput_payload_op1 = preRoundConstStage_input_payload_stateElement;
  assign preRoundConstStage_adderInput_payload_op2 = preRoundConstantMem_1_io_preConstant;
  assign preRoundConstStage_output_valid = preRoundConstStage_adderInst_io_output_valid;
  assign preRoundConstStage_output_payload_isFull = preRoundConstStage_addContextDelayed_isFull;
  assign preRoundConstStage_output_payload_fullRound = preRoundConstStage_addContextDelayed_fullRound;
  assign preRoundConstStage_output_payload_partialRound = preRoundConstStage_addContextDelayed_partialRound;
  assign preRoundConstStage_output_payload_stateIndex = preRoundConstStage_addContextDelayed_stateIndex;
  assign preRoundConstStage_output_payload_stateSize = preRoundConstStage_addContextDelayed_stateSize;
  assign preRoundConstStage_output_payload_stateID = preRoundConstStage_addContextDelayed_stateID;
  assign preRoundConstStage_output_payload_stateElements_0 = preRoundConstStage_addContextDelayed_stateElements_0;
  assign preRoundConstStage_output_payload_stateElements_1 = preRoundConstStage_addContextDelayed_stateElements_1;
  assign preRoundConstStage_output_payload_stateElements_2 = preRoundConstStage_addContextDelayed_stateElements_2;
  assign preRoundConstStage_output_payload_stateElements_3 = preRoundConstStage_addContextDelayed_stateElements_3;
  assign preRoundConstStage_output_payload_stateElements_4 = preRoundConstStage_addContextDelayed_stateElements_4;
  assign preRoundConstStage_output_payload_stateElements_5 = preRoundConstStage_addContextDelayed_stateElements_5;
  assign preRoundConstStage_output_payload_stateElements_6 = preRoundConstStage_addContextDelayed_stateElements_6;
  assign preRoundConstStage_output_payload_stateElements_7 = preRoundConstStage_addContextDelayed_stateElements_7;
  assign preRoundConstStage_output_payload_stateElements_8 = preRoundConstStage_addContextDelayed_stateElements_8;
  assign preRoundConstStage_output_payload_stateElements_9 = preRoundConstStage_addContextDelayed_stateElements_9;
  assign preRoundConstStage_output_payload_stateElements_10 = preRoundConstStage_addContextDelayed_stateElements_10;
  always @(*) begin
    preRoundConstStage_output_payload_stateElement = preRoundConstStage_addContextDelayed_stateElement;
    if(when_PoseidonTopLevel_l173) begin
      preRoundConstStage_output_payload_stateElement = preRoundConstStage_adderInst_io_output_payload_res;
    end
  end

  assign when_PoseidonTopLevel_l173 = (preRoundConstStage_addContextDelayed_fullRound == 3'b000);
  assign poseidonThread_1_io_output_toStream_valid = poseidonThread_1_io_output_valid;
  assign poseidonThread_1_io_output_toStream_payload_isFull = poseidonThread_1_io_output_payload_isFull;
  assign poseidonThread_1_io_output_toStream_payload_fullRound = poseidonThread_1_io_output_payload_fullRound;
  assign poseidonThread_1_io_output_toStream_payload_partialRound = poseidonThread_1_io_output_payload_partialRound;
  assign poseidonThread_1_io_output_toStream_payload_stateSize = poseidonThread_1_io_output_payload_stateSize;
  assign poseidonThread_1_io_output_toStream_payload_stateID = poseidonThread_1_io_output_payload_stateID;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_0 = poseidonThread_1_io_output_payload_stateElements_0;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_1 = poseidonThread_1_io_output_payload_stateElements_1;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_2 = poseidonThread_1_io_output_payload_stateElements_2;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_3 = poseidonThread_1_io_output_payload_stateElements_3;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_4 = poseidonThread_1_io_output_payload_stateElements_4;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_5 = poseidonThread_1_io_output_payload_stateElements_5;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_6 = poseidonThread_1_io_output_payload_stateElements_6;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_7 = poseidonThread_1_io_output_payload_stateElements_7;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_8 = poseidonThread_1_io_output_payload_stateElements_8;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_9 = poseidonThread_1_io_output_payload_stateElements_9;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_10 = poseidonThread_1_io_output_payload_stateElements_10;
  assign poseidonThread_1_io_output_toStream_payload_stateElements_11 = poseidonThread_1_io_output_payload_stateElements_11;
  assign poseidonThread_1_io_output_toStream_ready = demuxInst_io_input_ready;
  assign demuxInst_io_output0_ready = (! demuxInst_io_output0_rValid);
  assign demuxInst_io_output0_s2mPipe_valid = (demuxInst_io_output0_valid || demuxInst_io_output0_rValid);
  assign demuxInst_io_output0_s2mPipe_payload_isFull = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_isFull : demuxInst_io_output0_payload_isFull);
  assign demuxInst_io_output0_s2mPipe_payload_fullRound = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_fullRound : demuxInst_io_output0_payload_fullRound);
  assign demuxInst_io_output0_s2mPipe_payload_partialRound = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_partialRound : demuxInst_io_output0_payload_partialRound);
  assign demuxInst_io_output0_s2mPipe_payload_stateSize = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateSize : demuxInst_io_output0_payload_stateSize);
  assign demuxInst_io_output0_s2mPipe_payload_stateID = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateID : demuxInst_io_output0_payload_stateID);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_0 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_0 : demuxInst_io_output0_payload_stateElements_0);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_1 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_1 : demuxInst_io_output0_payload_stateElements_1);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_2 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_2 : demuxInst_io_output0_payload_stateElements_2);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_3 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_3 : demuxInst_io_output0_payload_stateElements_3);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_4 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_4 : demuxInst_io_output0_payload_stateElements_4);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_5 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_5 : demuxInst_io_output0_payload_stateElements_5);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_6 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_6 : demuxInst_io_output0_payload_stateElements_6);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_7 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_7 : demuxInst_io_output0_payload_stateElements_7);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_8 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_8 : demuxInst_io_output0_payload_stateElements_8);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_9 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_9 : demuxInst_io_output0_payload_stateElements_9);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_10 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_10 : demuxInst_io_output0_payload_stateElements_10);
  assign demuxInst_io_output0_s2mPipe_payload_stateElements_11 = (demuxInst_io_output0_rValid ? demuxInst_io_output0_rData_stateElements_11 : demuxInst_io_output0_payload_stateElements_11);
  always @(*) begin
    demuxInst_io_output0_s2mPipe_ready = loopback_ready;
    if(when_Stream_l342) begin
      demuxInst_io_output0_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! loopback_valid);
  assign loopback_valid = demuxInst_io_output0_s2mPipe_rValid;
  assign loopback_payload_isFull = demuxInst_io_output0_s2mPipe_rData_isFull;
  assign loopback_payload_fullRound = demuxInst_io_output0_s2mPipe_rData_fullRound;
  assign loopback_payload_partialRound = demuxInst_io_output0_s2mPipe_rData_partialRound;
  assign loopback_payload_stateSize = demuxInst_io_output0_s2mPipe_rData_stateSize;
  assign loopback_payload_stateID = demuxInst_io_output0_s2mPipe_rData_stateID;
  assign loopback_payload_stateElements_0 = demuxInst_io_output0_s2mPipe_rData_stateElements_0;
  assign loopback_payload_stateElements_1 = demuxInst_io_output0_s2mPipe_rData_stateElements_1;
  assign loopback_payload_stateElements_2 = demuxInst_io_output0_s2mPipe_rData_stateElements_2;
  assign loopback_payload_stateElements_3 = demuxInst_io_output0_s2mPipe_rData_stateElements_3;
  assign loopback_payload_stateElements_4 = demuxInst_io_output0_s2mPipe_rData_stateElements_4;
  assign loopback_payload_stateElements_5 = demuxInst_io_output0_s2mPipe_rData_stateElements_5;
  assign loopback_payload_stateElements_6 = demuxInst_io_output0_s2mPipe_rData_stateElements_6;
  assign loopback_payload_stateElements_7 = demuxInst_io_output0_s2mPipe_rData_stateElements_7;
  assign loopback_payload_stateElements_8 = demuxInst_io_output0_s2mPipe_rData_stateElements_8;
  assign loopback_payload_stateElements_9 = demuxInst_io_output0_s2mPipe_rData_stateElements_9;
  assign loopback_payload_stateElements_10 = demuxInst_io_output0_s2mPipe_rData_stateElements_10;
  assign loopback_payload_stateElements_11 = demuxInst_io_output0_s2mPipe_rData_stateElements_11;
  always @(*) begin
    demuxInst_io_output1_ready = demuxInst_io_output1_m2sPipe_ready;
    if(when_Stream_l342_1) begin
      demuxInst_io_output1_ready = 1'b1;
    end
  end

  assign when_Stream_l342_1 = (! demuxInst_io_output1_m2sPipe_valid);
  assign demuxInst_io_output1_m2sPipe_valid = demuxInst_io_output1_rValid;
  assign demuxInst_io_output1_m2sPipe_payload_stateID = demuxInst_io_output1_rData_stateID;
  assign demuxInst_io_output1_m2sPipe_payload_stateElement = demuxInst_io_output1_rData_stateElement;
  assign io_output_valid = demuxInst_io_output1_m2sPipe_valid;
  assign demuxInst_io_output1_m2sPipe_ready = io_output_ready;
  assign io_output_payload_stateID = demuxInst_io_output1_m2sPipe_payload_stateID;
  assign io_output_payload_stateElement = demuxInst_io_output1_m2sPipe_payload_stateElement;
  assign loopback_ready = bundleFifo_1_io_push_ready;
  assign loopbackBuffer_valid = bundleFifo_1_io_pop_valid;
  assign loopbackBuffer_payload_isFull = bundleFifo_1_io_pop_payload_isFull;
  assign loopbackBuffer_payload_fullRound = bundleFifo_1_io_pop_payload_fullRound;
  assign loopbackBuffer_payload_partialRound = bundleFifo_1_io_pop_payload_partialRound;
  assign loopbackBuffer_payload_stateSize = bundleFifo_1_io_pop_payload_stateSize;
  assign loopbackBuffer_payload_stateID = bundleFifo_1_io_pop_payload_stateID;
  assign loopbackBuffer_payload_stateElements_0 = bundleFifo_1_io_pop_payload_stateElements_0;
  assign loopbackBuffer_payload_stateElements_1 = bundleFifo_1_io_pop_payload_stateElements_1;
  assign loopbackBuffer_payload_stateElements_2 = bundleFifo_1_io_pop_payload_stateElements_2;
  assign loopbackBuffer_payload_stateElements_3 = bundleFifo_1_io_pop_payload_stateElements_3;
  assign loopbackBuffer_payload_stateElements_4 = bundleFifo_1_io_pop_payload_stateElements_4;
  assign loopbackBuffer_payload_stateElements_5 = bundleFifo_1_io_pop_payload_stateElements_5;
  assign loopbackBuffer_payload_stateElements_6 = bundleFifo_1_io_pop_payload_stateElements_6;
  assign loopbackBuffer_payload_stateElements_7 = bundleFifo_1_io_pop_payload_stateElements_7;
  assign loopbackBuffer_payload_stateElements_8 = bundleFifo_1_io_pop_payload_stateElements_8;
  assign loopbackBuffer_payload_stateElements_9 = bundleFifo_1_io_pop_payload_stateElements_9;
  assign loopbackBuffer_payload_stateElements_10 = bundleFifo_1_io_pop_payload_stateElements_10;
  assign loopbackBuffer_payload_stateElements_11 = bundleFifo_1_io_pop_payload_stateElements_11;
  always @(posedge clk) begin
    preRoundConstStage_input_payload_delay_1_isFull <= preRoundConstStage_input_payload_isFull;
    preRoundConstStage_input_payload_delay_1_fullRound <= preRoundConstStage_input_payload_fullRound;
    preRoundConstStage_input_payload_delay_1_partialRound <= preRoundConstStage_input_payload_partialRound;
    preRoundConstStage_input_payload_delay_1_stateIndex <= preRoundConstStage_input_payload_stateIndex;
    preRoundConstStage_input_payload_delay_1_stateSize <= preRoundConstStage_input_payload_stateSize;
    preRoundConstStage_input_payload_delay_1_stateID <= preRoundConstStage_input_payload_stateID;
    preRoundConstStage_input_payload_delay_1_stateElements_0 <= preRoundConstStage_input_payload_stateElements_0;
    preRoundConstStage_input_payload_delay_1_stateElements_1 <= preRoundConstStage_input_payload_stateElements_1;
    preRoundConstStage_input_payload_delay_1_stateElements_2 <= preRoundConstStage_input_payload_stateElements_2;
    preRoundConstStage_input_payload_delay_1_stateElements_3 <= preRoundConstStage_input_payload_stateElements_3;
    preRoundConstStage_input_payload_delay_1_stateElements_4 <= preRoundConstStage_input_payload_stateElements_4;
    preRoundConstStage_input_payload_delay_1_stateElements_5 <= preRoundConstStage_input_payload_stateElements_5;
    preRoundConstStage_input_payload_delay_1_stateElements_6 <= preRoundConstStage_input_payload_stateElements_6;
    preRoundConstStage_input_payload_delay_1_stateElements_7 <= preRoundConstStage_input_payload_stateElements_7;
    preRoundConstStage_input_payload_delay_1_stateElements_8 <= preRoundConstStage_input_payload_stateElements_8;
    preRoundConstStage_input_payload_delay_1_stateElements_9 <= preRoundConstStage_input_payload_stateElements_9;
    preRoundConstStage_input_payload_delay_1_stateElements_10 <= preRoundConstStage_input_payload_stateElements_10;
    preRoundConstStage_input_payload_delay_1_stateElement <= preRoundConstStage_input_payload_stateElement;
    preRoundConstStage_input_payload_delay_2_isFull <= preRoundConstStage_input_payload_delay_1_isFull;
    preRoundConstStage_input_payload_delay_2_fullRound <= preRoundConstStage_input_payload_delay_1_fullRound;
    preRoundConstStage_input_payload_delay_2_partialRound <= preRoundConstStage_input_payload_delay_1_partialRound;
    preRoundConstStage_input_payload_delay_2_stateIndex <= preRoundConstStage_input_payload_delay_1_stateIndex;
    preRoundConstStage_input_payload_delay_2_stateSize <= preRoundConstStage_input_payload_delay_1_stateSize;
    preRoundConstStage_input_payload_delay_2_stateID <= preRoundConstStage_input_payload_delay_1_stateID;
    preRoundConstStage_input_payload_delay_2_stateElements_0 <= preRoundConstStage_input_payload_delay_1_stateElements_0;
    preRoundConstStage_input_payload_delay_2_stateElements_1 <= preRoundConstStage_input_payload_delay_1_stateElements_1;
    preRoundConstStage_input_payload_delay_2_stateElements_2 <= preRoundConstStage_input_payload_delay_1_stateElements_2;
    preRoundConstStage_input_payload_delay_2_stateElements_3 <= preRoundConstStage_input_payload_delay_1_stateElements_3;
    preRoundConstStage_input_payload_delay_2_stateElements_4 <= preRoundConstStage_input_payload_delay_1_stateElements_4;
    preRoundConstStage_input_payload_delay_2_stateElements_5 <= preRoundConstStage_input_payload_delay_1_stateElements_5;
    preRoundConstStage_input_payload_delay_2_stateElements_6 <= preRoundConstStage_input_payload_delay_1_stateElements_6;
    preRoundConstStage_input_payload_delay_2_stateElements_7 <= preRoundConstStage_input_payload_delay_1_stateElements_7;
    preRoundConstStage_input_payload_delay_2_stateElements_8 <= preRoundConstStage_input_payload_delay_1_stateElements_8;
    preRoundConstStage_input_payload_delay_2_stateElements_9 <= preRoundConstStage_input_payload_delay_1_stateElements_9;
    preRoundConstStage_input_payload_delay_2_stateElements_10 <= preRoundConstStage_input_payload_delay_1_stateElements_10;
    preRoundConstStage_input_payload_delay_2_stateElement <= preRoundConstStage_input_payload_delay_1_stateElement;
    preRoundConstStage_input_payload_delay_3_isFull <= preRoundConstStage_input_payload_delay_2_isFull;
    preRoundConstStage_input_payload_delay_3_fullRound <= preRoundConstStage_input_payload_delay_2_fullRound;
    preRoundConstStage_input_payload_delay_3_partialRound <= preRoundConstStage_input_payload_delay_2_partialRound;
    preRoundConstStage_input_payload_delay_3_stateIndex <= preRoundConstStage_input_payload_delay_2_stateIndex;
    preRoundConstStage_input_payload_delay_3_stateSize <= preRoundConstStage_input_payload_delay_2_stateSize;
    preRoundConstStage_input_payload_delay_3_stateID <= preRoundConstStage_input_payload_delay_2_stateID;
    preRoundConstStage_input_payload_delay_3_stateElements_0 <= preRoundConstStage_input_payload_delay_2_stateElements_0;
    preRoundConstStage_input_payload_delay_3_stateElements_1 <= preRoundConstStage_input_payload_delay_2_stateElements_1;
    preRoundConstStage_input_payload_delay_3_stateElements_2 <= preRoundConstStage_input_payload_delay_2_stateElements_2;
    preRoundConstStage_input_payload_delay_3_stateElements_3 <= preRoundConstStage_input_payload_delay_2_stateElements_3;
    preRoundConstStage_input_payload_delay_3_stateElements_4 <= preRoundConstStage_input_payload_delay_2_stateElements_4;
    preRoundConstStage_input_payload_delay_3_stateElements_5 <= preRoundConstStage_input_payload_delay_2_stateElements_5;
    preRoundConstStage_input_payload_delay_3_stateElements_6 <= preRoundConstStage_input_payload_delay_2_stateElements_6;
    preRoundConstStage_input_payload_delay_3_stateElements_7 <= preRoundConstStage_input_payload_delay_2_stateElements_7;
    preRoundConstStage_input_payload_delay_3_stateElements_8 <= preRoundConstStage_input_payload_delay_2_stateElements_8;
    preRoundConstStage_input_payload_delay_3_stateElements_9 <= preRoundConstStage_input_payload_delay_2_stateElements_9;
    preRoundConstStage_input_payload_delay_3_stateElements_10 <= preRoundConstStage_input_payload_delay_2_stateElements_10;
    preRoundConstStage_input_payload_delay_3_stateElement <= preRoundConstStage_input_payload_delay_2_stateElement;
    preRoundConstStage_input_payload_delay_4_isFull <= preRoundConstStage_input_payload_delay_3_isFull;
    preRoundConstStage_input_payload_delay_4_fullRound <= preRoundConstStage_input_payload_delay_3_fullRound;
    preRoundConstStage_input_payload_delay_4_partialRound <= preRoundConstStage_input_payload_delay_3_partialRound;
    preRoundConstStage_input_payload_delay_4_stateIndex <= preRoundConstStage_input_payload_delay_3_stateIndex;
    preRoundConstStage_input_payload_delay_4_stateSize <= preRoundConstStage_input_payload_delay_3_stateSize;
    preRoundConstStage_input_payload_delay_4_stateID <= preRoundConstStage_input_payload_delay_3_stateID;
    preRoundConstStage_input_payload_delay_4_stateElements_0 <= preRoundConstStage_input_payload_delay_3_stateElements_0;
    preRoundConstStage_input_payload_delay_4_stateElements_1 <= preRoundConstStage_input_payload_delay_3_stateElements_1;
    preRoundConstStage_input_payload_delay_4_stateElements_2 <= preRoundConstStage_input_payload_delay_3_stateElements_2;
    preRoundConstStage_input_payload_delay_4_stateElements_3 <= preRoundConstStage_input_payload_delay_3_stateElements_3;
    preRoundConstStage_input_payload_delay_4_stateElements_4 <= preRoundConstStage_input_payload_delay_3_stateElements_4;
    preRoundConstStage_input_payload_delay_4_stateElements_5 <= preRoundConstStage_input_payload_delay_3_stateElements_5;
    preRoundConstStage_input_payload_delay_4_stateElements_6 <= preRoundConstStage_input_payload_delay_3_stateElements_6;
    preRoundConstStage_input_payload_delay_4_stateElements_7 <= preRoundConstStage_input_payload_delay_3_stateElements_7;
    preRoundConstStage_input_payload_delay_4_stateElements_8 <= preRoundConstStage_input_payload_delay_3_stateElements_8;
    preRoundConstStage_input_payload_delay_4_stateElements_9 <= preRoundConstStage_input_payload_delay_3_stateElements_9;
    preRoundConstStage_input_payload_delay_4_stateElements_10 <= preRoundConstStage_input_payload_delay_3_stateElements_10;
    preRoundConstStage_input_payload_delay_4_stateElement <= preRoundConstStage_input_payload_delay_3_stateElement;
    preRoundConstStage_input_payload_delay_5_isFull <= preRoundConstStage_input_payload_delay_4_isFull;
    preRoundConstStage_input_payload_delay_5_fullRound <= preRoundConstStage_input_payload_delay_4_fullRound;
    preRoundConstStage_input_payload_delay_5_partialRound <= preRoundConstStage_input_payload_delay_4_partialRound;
    preRoundConstStage_input_payload_delay_5_stateIndex <= preRoundConstStage_input_payload_delay_4_stateIndex;
    preRoundConstStage_input_payload_delay_5_stateSize <= preRoundConstStage_input_payload_delay_4_stateSize;
    preRoundConstStage_input_payload_delay_5_stateID <= preRoundConstStage_input_payload_delay_4_stateID;
    preRoundConstStage_input_payload_delay_5_stateElements_0 <= preRoundConstStage_input_payload_delay_4_stateElements_0;
    preRoundConstStage_input_payload_delay_5_stateElements_1 <= preRoundConstStage_input_payload_delay_4_stateElements_1;
    preRoundConstStage_input_payload_delay_5_stateElements_2 <= preRoundConstStage_input_payload_delay_4_stateElements_2;
    preRoundConstStage_input_payload_delay_5_stateElements_3 <= preRoundConstStage_input_payload_delay_4_stateElements_3;
    preRoundConstStage_input_payload_delay_5_stateElements_4 <= preRoundConstStage_input_payload_delay_4_stateElements_4;
    preRoundConstStage_input_payload_delay_5_stateElements_5 <= preRoundConstStage_input_payload_delay_4_stateElements_5;
    preRoundConstStage_input_payload_delay_5_stateElements_6 <= preRoundConstStage_input_payload_delay_4_stateElements_6;
    preRoundConstStage_input_payload_delay_5_stateElements_7 <= preRoundConstStage_input_payload_delay_4_stateElements_7;
    preRoundConstStage_input_payload_delay_5_stateElements_8 <= preRoundConstStage_input_payload_delay_4_stateElements_8;
    preRoundConstStage_input_payload_delay_5_stateElements_9 <= preRoundConstStage_input_payload_delay_4_stateElements_9;
    preRoundConstStage_input_payload_delay_5_stateElements_10 <= preRoundConstStage_input_payload_delay_4_stateElements_10;
    preRoundConstStage_input_payload_delay_5_stateElement <= preRoundConstStage_input_payload_delay_4_stateElement;
    preRoundConstStage_input_payload_delay_6_isFull <= preRoundConstStage_input_payload_delay_5_isFull;
    preRoundConstStage_input_payload_delay_6_fullRound <= preRoundConstStage_input_payload_delay_5_fullRound;
    preRoundConstStage_input_payload_delay_6_partialRound <= preRoundConstStage_input_payload_delay_5_partialRound;
    preRoundConstStage_input_payload_delay_6_stateIndex <= preRoundConstStage_input_payload_delay_5_stateIndex;
    preRoundConstStage_input_payload_delay_6_stateSize <= preRoundConstStage_input_payload_delay_5_stateSize;
    preRoundConstStage_input_payload_delay_6_stateID <= preRoundConstStage_input_payload_delay_5_stateID;
    preRoundConstStage_input_payload_delay_6_stateElements_0 <= preRoundConstStage_input_payload_delay_5_stateElements_0;
    preRoundConstStage_input_payload_delay_6_stateElements_1 <= preRoundConstStage_input_payload_delay_5_stateElements_1;
    preRoundConstStage_input_payload_delay_6_stateElements_2 <= preRoundConstStage_input_payload_delay_5_stateElements_2;
    preRoundConstStage_input_payload_delay_6_stateElements_3 <= preRoundConstStage_input_payload_delay_5_stateElements_3;
    preRoundConstStage_input_payload_delay_6_stateElements_4 <= preRoundConstStage_input_payload_delay_5_stateElements_4;
    preRoundConstStage_input_payload_delay_6_stateElements_5 <= preRoundConstStage_input_payload_delay_5_stateElements_5;
    preRoundConstStage_input_payload_delay_6_stateElements_6 <= preRoundConstStage_input_payload_delay_5_stateElements_6;
    preRoundConstStage_input_payload_delay_6_stateElements_7 <= preRoundConstStage_input_payload_delay_5_stateElements_7;
    preRoundConstStage_input_payload_delay_6_stateElements_8 <= preRoundConstStage_input_payload_delay_5_stateElements_8;
    preRoundConstStage_input_payload_delay_6_stateElements_9 <= preRoundConstStage_input_payload_delay_5_stateElements_9;
    preRoundConstStage_input_payload_delay_6_stateElements_10 <= preRoundConstStage_input_payload_delay_5_stateElements_10;
    preRoundConstStage_input_payload_delay_6_stateElement <= preRoundConstStage_input_payload_delay_5_stateElement;
    preRoundConstStage_input_payload_delay_7_isFull <= preRoundConstStage_input_payload_delay_6_isFull;
    preRoundConstStage_input_payload_delay_7_fullRound <= preRoundConstStage_input_payload_delay_6_fullRound;
    preRoundConstStage_input_payload_delay_7_partialRound <= preRoundConstStage_input_payload_delay_6_partialRound;
    preRoundConstStage_input_payload_delay_7_stateIndex <= preRoundConstStage_input_payload_delay_6_stateIndex;
    preRoundConstStage_input_payload_delay_7_stateSize <= preRoundConstStage_input_payload_delay_6_stateSize;
    preRoundConstStage_input_payload_delay_7_stateID <= preRoundConstStage_input_payload_delay_6_stateID;
    preRoundConstStage_input_payload_delay_7_stateElements_0 <= preRoundConstStage_input_payload_delay_6_stateElements_0;
    preRoundConstStage_input_payload_delay_7_stateElements_1 <= preRoundConstStage_input_payload_delay_6_stateElements_1;
    preRoundConstStage_input_payload_delay_7_stateElements_2 <= preRoundConstStage_input_payload_delay_6_stateElements_2;
    preRoundConstStage_input_payload_delay_7_stateElements_3 <= preRoundConstStage_input_payload_delay_6_stateElements_3;
    preRoundConstStage_input_payload_delay_7_stateElements_4 <= preRoundConstStage_input_payload_delay_6_stateElements_4;
    preRoundConstStage_input_payload_delay_7_stateElements_5 <= preRoundConstStage_input_payload_delay_6_stateElements_5;
    preRoundConstStage_input_payload_delay_7_stateElements_6 <= preRoundConstStage_input_payload_delay_6_stateElements_6;
    preRoundConstStage_input_payload_delay_7_stateElements_7 <= preRoundConstStage_input_payload_delay_6_stateElements_7;
    preRoundConstStage_input_payload_delay_7_stateElements_8 <= preRoundConstStage_input_payload_delay_6_stateElements_8;
    preRoundConstStage_input_payload_delay_7_stateElements_9 <= preRoundConstStage_input_payload_delay_6_stateElements_9;
    preRoundConstStage_input_payload_delay_7_stateElements_10 <= preRoundConstStage_input_payload_delay_6_stateElements_10;
    preRoundConstStage_input_payload_delay_7_stateElement <= preRoundConstStage_input_payload_delay_6_stateElement;
    preRoundConstStage_input_payload_delay_8_isFull <= preRoundConstStage_input_payload_delay_7_isFull;
    preRoundConstStage_input_payload_delay_8_fullRound <= preRoundConstStage_input_payload_delay_7_fullRound;
    preRoundConstStage_input_payload_delay_8_partialRound <= preRoundConstStage_input_payload_delay_7_partialRound;
    preRoundConstStage_input_payload_delay_8_stateIndex <= preRoundConstStage_input_payload_delay_7_stateIndex;
    preRoundConstStage_input_payload_delay_8_stateSize <= preRoundConstStage_input_payload_delay_7_stateSize;
    preRoundConstStage_input_payload_delay_8_stateID <= preRoundConstStage_input_payload_delay_7_stateID;
    preRoundConstStage_input_payload_delay_8_stateElements_0 <= preRoundConstStage_input_payload_delay_7_stateElements_0;
    preRoundConstStage_input_payload_delay_8_stateElements_1 <= preRoundConstStage_input_payload_delay_7_stateElements_1;
    preRoundConstStage_input_payload_delay_8_stateElements_2 <= preRoundConstStage_input_payload_delay_7_stateElements_2;
    preRoundConstStage_input_payload_delay_8_stateElements_3 <= preRoundConstStage_input_payload_delay_7_stateElements_3;
    preRoundConstStage_input_payload_delay_8_stateElements_4 <= preRoundConstStage_input_payload_delay_7_stateElements_4;
    preRoundConstStage_input_payload_delay_8_stateElements_5 <= preRoundConstStage_input_payload_delay_7_stateElements_5;
    preRoundConstStage_input_payload_delay_8_stateElements_6 <= preRoundConstStage_input_payload_delay_7_stateElements_6;
    preRoundConstStage_input_payload_delay_8_stateElements_7 <= preRoundConstStage_input_payload_delay_7_stateElements_7;
    preRoundConstStage_input_payload_delay_8_stateElements_8 <= preRoundConstStage_input_payload_delay_7_stateElements_8;
    preRoundConstStage_input_payload_delay_8_stateElements_9 <= preRoundConstStage_input_payload_delay_7_stateElements_9;
    preRoundConstStage_input_payload_delay_8_stateElements_10 <= preRoundConstStage_input_payload_delay_7_stateElements_10;
    preRoundConstStage_input_payload_delay_8_stateElement <= preRoundConstStage_input_payload_delay_7_stateElement;
    preRoundConstStage_input_payload_delay_9_isFull <= preRoundConstStage_input_payload_delay_8_isFull;
    preRoundConstStage_input_payload_delay_9_fullRound <= preRoundConstStage_input_payload_delay_8_fullRound;
    preRoundConstStage_input_payload_delay_9_partialRound <= preRoundConstStage_input_payload_delay_8_partialRound;
    preRoundConstStage_input_payload_delay_9_stateIndex <= preRoundConstStage_input_payload_delay_8_stateIndex;
    preRoundConstStage_input_payload_delay_9_stateSize <= preRoundConstStage_input_payload_delay_8_stateSize;
    preRoundConstStage_input_payload_delay_9_stateID <= preRoundConstStage_input_payload_delay_8_stateID;
    preRoundConstStage_input_payload_delay_9_stateElements_0 <= preRoundConstStage_input_payload_delay_8_stateElements_0;
    preRoundConstStage_input_payload_delay_9_stateElements_1 <= preRoundConstStage_input_payload_delay_8_stateElements_1;
    preRoundConstStage_input_payload_delay_9_stateElements_2 <= preRoundConstStage_input_payload_delay_8_stateElements_2;
    preRoundConstStage_input_payload_delay_9_stateElements_3 <= preRoundConstStage_input_payload_delay_8_stateElements_3;
    preRoundConstStage_input_payload_delay_9_stateElements_4 <= preRoundConstStage_input_payload_delay_8_stateElements_4;
    preRoundConstStage_input_payload_delay_9_stateElements_5 <= preRoundConstStage_input_payload_delay_8_stateElements_5;
    preRoundConstStage_input_payload_delay_9_stateElements_6 <= preRoundConstStage_input_payload_delay_8_stateElements_6;
    preRoundConstStage_input_payload_delay_9_stateElements_7 <= preRoundConstStage_input_payload_delay_8_stateElements_7;
    preRoundConstStage_input_payload_delay_9_stateElements_8 <= preRoundConstStage_input_payload_delay_8_stateElements_8;
    preRoundConstStage_input_payload_delay_9_stateElements_9 <= preRoundConstStage_input_payload_delay_8_stateElements_9;
    preRoundConstStage_input_payload_delay_9_stateElements_10 <= preRoundConstStage_input_payload_delay_8_stateElements_10;
    preRoundConstStage_input_payload_delay_9_stateElement <= preRoundConstStage_input_payload_delay_8_stateElement;
    preRoundConstStage_input_payload_delay_10_isFull <= preRoundConstStage_input_payload_delay_9_isFull;
    preRoundConstStage_input_payload_delay_10_fullRound <= preRoundConstStage_input_payload_delay_9_fullRound;
    preRoundConstStage_input_payload_delay_10_partialRound <= preRoundConstStage_input_payload_delay_9_partialRound;
    preRoundConstStage_input_payload_delay_10_stateIndex <= preRoundConstStage_input_payload_delay_9_stateIndex;
    preRoundConstStage_input_payload_delay_10_stateSize <= preRoundConstStage_input_payload_delay_9_stateSize;
    preRoundConstStage_input_payload_delay_10_stateID <= preRoundConstStage_input_payload_delay_9_stateID;
    preRoundConstStage_input_payload_delay_10_stateElements_0 <= preRoundConstStage_input_payload_delay_9_stateElements_0;
    preRoundConstStage_input_payload_delay_10_stateElements_1 <= preRoundConstStage_input_payload_delay_9_stateElements_1;
    preRoundConstStage_input_payload_delay_10_stateElements_2 <= preRoundConstStage_input_payload_delay_9_stateElements_2;
    preRoundConstStage_input_payload_delay_10_stateElements_3 <= preRoundConstStage_input_payload_delay_9_stateElements_3;
    preRoundConstStage_input_payload_delay_10_stateElements_4 <= preRoundConstStage_input_payload_delay_9_stateElements_4;
    preRoundConstStage_input_payload_delay_10_stateElements_5 <= preRoundConstStage_input_payload_delay_9_stateElements_5;
    preRoundConstStage_input_payload_delay_10_stateElements_6 <= preRoundConstStage_input_payload_delay_9_stateElements_6;
    preRoundConstStage_input_payload_delay_10_stateElements_7 <= preRoundConstStage_input_payload_delay_9_stateElements_7;
    preRoundConstStage_input_payload_delay_10_stateElements_8 <= preRoundConstStage_input_payload_delay_9_stateElements_8;
    preRoundConstStage_input_payload_delay_10_stateElements_9 <= preRoundConstStage_input_payload_delay_9_stateElements_9;
    preRoundConstStage_input_payload_delay_10_stateElements_10 <= preRoundConstStage_input_payload_delay_9_stateElements_10;
    preRoundConstStage_input_payload_delay_10_stateElement <= preRoundConstStage_input_payload_delay_9_stateElement;
    preRoundConstStage_input_payload_delay_11_isFull <= preRoundConstStage_input_payload_delay_10_isFull;
    preRoundConstStage_input_payload_delay_11_fullRound <= preRoundConstStage_input_payload_delay_10_fullRound;
    preRoundConstStage_input_payload_delay_11_partialRound <= preRoundConstStage_input_payload_delay_10_partialRound;
    preRoundConstStage_input_payload_delay_11_stateIndex <= preRoundConstStage_input_payload_delay_10_stateIndex;
    preRoundConstStage_input_payload_delay_11_stateSize <= preRoundConstStage_input_payload_delay_10_stateSize;
    preRoundConstStage_input_payload_delay_11_stateID <= preRoundConstStage_input_payload_delay_10_stateID;
    preRoundConstStage_input_payload_delay_11_stateElements_0 <= preRoundConstStage_input_payload_delay_10_stateElements_0;
    preRoundConstStage_input_payload_delay_11_stateElements_1 <= preRoundConstStage_input_payload_delay_10_stateElements_1;
    preRoundConstStage_input_payload_delay_11_stateElements_2 <= preRoundConstStage_input_payload_delay_10_stateElements_2;
    preRoundConstStage_input_payload_delay_11_stateElements_3 <= preRoundConstStage_input_payload_delay_10_stateElements_3;
    preRoundConstStage_input_payload_delay_11_stateElements_4 <= preRoundConstStage_input_payload_delay_10_stateElements_4;
    preRoundConstStage_input_payload_delay_11_stateElements_5 <= preRoundConstStage_input_payload_delay_10_stateElements_5;
    preRoundConstStage_input_payload_delay_11_stateElements_6 <= preRoundConstStage_input_payload_delay_10_stateElements_6;
    preRoundConstStage_input_payload_delay_11_stateElements_7 <= preRoundConstStage_input_payload_delay_10_stateElements_7;
    preRoundConstStage_input_payload_delay_11_stateElements_8 <= preRoundConstStage_input_payload_delay_10_stateElements_8;
    preRoundConstStage_input_payload_delay_11_stateElements_9 <= preRoundConstStage_input_payload_delay_10_stateElements_9;
    preRoundConstStage_input_payload_delay_11_stateElements_10 <= preRoundConstStage_input_payload_delay_10_stateElements_10;
    preRoundConstStage_input_payload_delay_11_stateElement <= preRoundConstStage_input_payload_delay_10_stateElement;
    preRoundConstStage_input_payload_delay_12_isFull <= preRoundConstStage_input_payload_delay_11_isFull;
    preRoundConstStage_input_payload_delay_12_fullRound <= preRoundConstStage_input_payload_delay_11_fullRound;
    preRoundConstStage_input_payload_delay_12_partialRound <= preRoundConstStage_input_payload_delay_11_partialRound;
    preRoundConstStage_input_payload_delay_12_stateIndex <= preRoundConstStage_input_payload_delay_11_stateIndex;
    preRoundConstStage_input_payload_delay_12_stateSize <= preRoundConstStage_input_payload_delay_11_stateSize;
    preRoundConstStage_input_payload_delay_12_stateID <= preRoundConstStage_input_payload_delay_11_stateID;
    preRoundConstStage_input_payload_delay_12_stateElements_0 <= preRoundConstStage_input_payload_delay_11_stateElements_0;
    preRoundConstStage_input_payload_delay_12_stateElements_1 <= preRoundConstStage_input_payload_delay_11_stateElements_1;
    preRoundConstStage_input_payload_delay_12_stateElements_2 <= preRoundConstStage_input_payload_delay_11_stateElements_2;
    preRoundConstStage_input_payload_delay_12_stateElements_3 <= preRoundConstStage_input_payload_delay_11_stateElements_3;
    preRoundConstStage_input_payload_delay_12_stateElements_4 <= preRoundConstStage_input_payload_delay_11_stateElements_4;
    preRoundConstStage_input_payload_delay_12_stateElements_5 <= preRoundConstStage_input_payload_delay_11_stateElements_5;
    preRoundConstStage_input_payload_delay_12_stateElements_6 <= preRoundConstStage_input_payload_delay_11_stateElements_6;
    preRoundConstStage_input_payload_delay_12_stateElements_7 <= preRoundConstStage_input_payload_delay_11_stateElements_7;
    preRoundConstStage_input_payload_delay_12_stateElements_8 <= preRoundConstStage_input_payload_delay_11_stateElements_8;
    preRoundConstStage_input_payload_delay_12_stateElements_9 <= preRoundConstStage_input_payload_delay_11_stateElements_9;
    preRoundConstStage_input_payload_delay_12_stateElements_10 <= preRoundConstStage_input_payload_delay_11_stateElements_10;
    preRoundConstStage_input_payload_delay_12_stateElement <= preRoundConstStage_input_payload_delay_11_stateElement;
    preRoundConstStage_input_payload_delay_13_isFull <= preRoundConstStage_input_payload_delay_12_isFull;
    preRoundConstStage_input_payload_delay_13_fullRound <= preRoundConstStage_input_payload_delay_12_fullRound;
    preRoundConstStage_input_payload_delay_13_partialRound <= preRoundConstStage_input_payload_delay_12_partialRound;
    preRoundConstStage_input_payload_delay_13_stateIndex <= preRoundConstStage_input_payload_delay_12_stateIndex;
    preRoundConstStage_input_payload_delay_13_stateSize <= preRoundConstStage_input_payload_delay_12_stateSize;
    preRoundConstStage_input_payload_delay_13_stateID <= preRoundConstStage_input_payload_delay_12_stateID;
    preRoundConstStage_input_payload_delay_13_stateElements_0 <= preRoundConstStage_input_payload_delay_12_stateElements_0;
    preRoundConstStage_input_payload_delay_13_stateElements_1 <= preRoundConstStage_input_payload_delay_12_stateElements_1;
    preRoundConstStage_input_payload_delay_13_stateElements_2 <= preRoundConstStage_input_payload_delay_12_stateElements_2;
    preRoundConstStage_input_payload_delay_13_stateElements_3 <= preRoundConstStage_input_payload_delay_12_stateElements_3;
    preRoundConstStage_input_payload_delay_13_stateElements_4 <= preRoundConstStage_input_payload_delay_12_stateElements_4;
    preRoundConstStage_input_payload_delay_13_stateElements_5 <= preRoundConstStage_input_payload_delay_12_stateElements_5;
    preRoundConstStage_input_payload_delay_13_stateElements_6 <= preRoundConstStage_input_payload_delay_12_stateElements_6;
    preRoundConstStage_input_payload_delay_13_stateElements_7 <= preRoundConstStage_input_payload_delay_12_stateElements_7;
    preRoundConstStage_input_payload_delay_13_stateElements_8 <= preRoundConstStage_input_payload_delay_12_stateElements_8;
    preRoundConstStage_input_payload_delay_13_stateElements_9 <= preRoundConstStage_input_payload_delay_12_stateElements_9;
    preRoundConstStage_input_payload_delay_13_stateElements_10 <= preRoundConstStage_input_payload_delay_12_stateElements_10;
    preRoundConstStage_input_payload_delay_13_stateElement <= preRoundConstStage_input_payload_delay_12_stateElement;
    preRoundConstStage_input_payload_delay_14_isFull <= preRoundConstStage_input_payload_delay_13_isFull;
    preRoundConstStage_input_payload_delay_14_fullRound <= preRoundConstStage_input_payload_delay_13_fullRound;
    preRoundConstStage_input_payload_delay_14_partialRound <= preRoundConstStage_input_payload_delay_13_partialRound;
    preRoundConstStage_input_payload_delay_14_stateIndex <= preRoundConstStage_input_payload_delay_13_stateIndex;
    preRoundConstStage_input_payload_delay_14_stateSize <= preRoundConstStage_input_payload_delay_13_stateSize;
    preRoundConstStage_input_payload_delay_14_stateID <= preRoundConstStage_input_payload_delay_13_stateID;
    preRoundConstStage_input_payload_delay_14_stateElements_0 <= preRoundConstStage_input_payload_delay_13_stateElements_0;
    preRoundConstStage_input_payload_delay_14_stateElements_1 <= preRoundConstStage_input_payload_delay_13_stateElements_1;
    preRoundConstStage_input_payload_delay_14_stateElements_2 <= preRoundConstStage_input_payload_delay_13_stateElements_2;
    preRoundConstStage_input_payload_delay_14_stateElements_3 <= preRoundConstStage_input_payload_delay_13_stateElements_3;
    preRoundConstStage_input_payload_delay_14_stateElements_4 <= preRoundConstStage_input_payload_delay_13_stateElements_4;
    preRoundConstStage_input_payload_delay_14_stateElements_5 <= preRoundConstStage_input_payload_delay_13_stateElements_5;
    preRoundConstStage_input_payload_delay_14_stateElements_6 <= preRoundConstStage_input_payload_delay_13_stateElements_6;
    preRoundConstStage_input_payload_delay_14_stateElements_7 <= preRoundConstStage_input_payload_delay_13_stateElements_7;
    preRoundConstStage_input_payload_delay_14_stateElements_8 <= preRoundConstStage_input_payload_delay_13_stateElements_8;
    preRoundConstStage_input_payload_delay_14_stateElements_9 <= preRoundConstStage_input_payload_delay_13_stateElements_9;
    preRoundConstStage_input_payload_delay_14_stateElements_10 <= preRoundConstStage_input_payload_delay_13_stateElements_10;
    preRoundConstStage_input_payload_delay_14_stateElement <= preRoundConstStage_input_payload_delay_13_stateElement;
    preRoundConstStage_input_payload_delay_15_isFull <= preRoundConstStage_input_payload_delay_14_isFull;
    preRoundConstStage_input_payload_delay_15_fullRound <= preRoundConstStage_input_payload_delay_14_fullRound;
    preRoundConstStage_input_payload_delay_15_partialRound <= preRoundConstStage_input_payload_delay_14_partialRound;
    preRoundConstStage_input_payload_delay_15_stateIndex <= preRoundConstStage_input_payload_delay_14_stateIndex;
    preRoundConstStage_input_payload_delay_15_stateSize <= preRoundConstStage_input_payload_delay_14_stateSize;
    preRoundConstStage_input_payload_delay_15_stateID <= preRoundConstStage_input_payload_delay_14_stateID;
    preRoundConstStage_input_payload_delay_15_stateElements_0 <= preRoundConstStage_input_payload_delay_14_stateElements_0;
    preRoundConstStage_input_payload_delay_15_stateElements_1 <= preRoundConstStage_input_payload_delay_14_stateElements_1;
    preRoundConstStage_input_payload_delay_15_stateElements_2 <= preRoundConstStage_input_payload_delay_14_stateElements_2;
    preRoundConstStage_input_payload_delay_15_stateElements_3 <= preRoundConstStage_input_payload_delay_14_stateElements_3;
    preRoundConstStage_input_payload_delay_15_stateElements_4 <= preRoundConstStage_input_payload_delay_14_stateElements_4;
    preRoundConstStage_input_payload_delay_15_stateElements_5 <= preRoundConstStage_input_payload_delay_14_stateElements_5;
    preRoundConstStage_input_payload_delay_15_stateElements_6 <= preRoundConstStage_input_payload_delay_14_stateElements_6;
    preRoundConstStage_input_payload_delay_15_stateElements_7 <= preRoundConstStage_input_payload_delay_14_stateElements_7;
    preRoundConstStage_input_payload_delay_15_stateElements_8 <= preRoundConstStage_input_payload_delay_14_stateElements_8;
    preRoundConstStage_input_payload_delay_15_stateElements_9 <= preRoundConstStage_input_payload_delay_14_stateElements_9;
    preRoundConstStage_input_payload_delay_15_stateElements_10 <= preRoundConstStage_input_payload_delay_14_stateElements_10;
    preRoundConstStage_input_payload_delay_15_stateElement <= preRoundConstStage_input_payload_delay_14_stateElement;
    preRoundConstStage_input_payload_delay_16_isFull <= preRoundConstStage_input_payload_delay_15_isFull;
    preRoundConstStage_input_payload_delay_16_fullRound <= preRoundConstStage_input_payload_delay_15_fullRound;
    preRoundConstStage_input_payload_delay_16_partialRound <= preRoundConstStage_input_payload_delay_15_partialRound;
    preRoundConstStage_input_payload_delay_16_stateIndex <= preRoundConstStage_input_payload_delay_15_stateIndex;
    preRoundConstStage_input_payload_delay_16_stateSize <= preRoundConstStage_input_payload_delay_15_stateSize;
    preRoundConstStage_input_payload_delay_16_stateID <= preRoundConstStage_input_payload_delay_15_stateID;
    preRoundConstStage_input_payload_delay_16_stateElements_0 <= preRoundConstStage_input_payload_delay_15_stateElements_0;
    preRoundConstStage_input_payload_delay_16_stateElements_1 <= preRoundConstStage_input_payload_delay_15_stateElements_1;
    preRoundConstStage_input_payload_delay_16_stateElements_2 <= preRoundConstStage_input_payload_delay_15_stateElements_2;
    preRoundConstStage_input_payload_delay_16_stateElements_3 <= preRoundConstStage_input_payload_delay_15_stateElements_3;
    preRoundConstStage_input_payload_delay_16_stateElements_4 <= preRoundConstStage_input_payload_delay_15_stateElements_4;
    preRoundConstStage_input_payload_delay_16_stateElements_5 <= preRoundConstStage_input_payload_delay_15_stateElements_5;
    preRoundConstStage_input_payload_delay_16_stateElements_6 <= preRoundConstStage_input_payload_delay_15_stateElements_6;
    preRoundConstStage_input_payload_delay_16_stateElements_7 <= preRoundConstStage_input_payload_delay_15_stateElements_7;
    preRoundConstStage_input_payload_delay_16_stateElements_8 <= preRoundConstStage_input_payload_delay_15_stateElements_8;
    preRoundConstStage_input_payload_delay_16_stateElements_9 <= preRoundConstStage_input_payload_delay_15_stateElements_9;
    preRoundConstStage_input_payload_delay_16_stateElements_10 <= preRoundConstStage_input_payload_delay_15_stateElements_10;
    preRoundConstStage_input_payload_delay_16_stateElement <= preRoundConstStage_input_payload_delay_15_stateElement;
    preRoundConstStage_addContextDelayed_isFull <= preRoundConstStage_input_payload_delay_16_isFull;
    preRoundConstStage_addContextDelayed_fullRound <= preRoundConstStage_input_payload_delay_16_fullRound;
    preRoundConstStage_addContextDelayed_partialRound <= preRoundConstStage_input_payload_delay_16_partialRound;
    preRoundConstStage_addContextDelayed_stateIndex <= preRoundConstStage_input_payload_delay_16_stateIndex;
    preRoundConstStage_addContextDelayed_stateSize <= preRoundConstStage_input_payload_delay_16_stateSize;
    preRoundConstStage_addContextDelayed_stateID <= preRoundConstStage_input_payload_delay_16_stateID;
    preRoundConstStage_addContextDelayed_stateElements_0 <= preRoundConstStage_input_payload_delay_16_stateElements_0;
    preRoundConstStage_addContextDelayed_stateElements_1 <= preRoundConstStage_input_payload_delay_16_stateElements_1;
    preRoundConstStage_addContextDelayed_stateElements_2 <= preRoundConstStage_input_payload_delay_16_stateElements_2;
    preRoundConstStage_addContextDelayed_stateElements_3 <= preRoundConstStage_input_payload_delay_16_stateElements_3;
    preRoundConstStage_addContextDelayed_stateElements_4 <= preRoundConstStage_input_payload_delay_16_stateElements_4;
    preRoundConstStage_addContextDelayed_stateElements_5 <= preRoundConstStage_input_payload_delay_16_stateElements_5;
    preRoundConstStage_addContextDelayed_stateElements_6 <= preRoundConstStage_input_payload_delay_16_stateElements_6;
    preRoundConstStage_addContextDelayed_stateElements_7 <= preRoundConstStage_input_payload_delay_16_stateElements_7;
    preRoundConstStage_addContextDelayed_stateElements_8 <= preRoundConstStage_input_payload_delay_16_stateElements_8;
    preRoundConstStage_addContextDelayed_stateElements_9 <= preRoundConstStage_input_payload_delay_16_stateElements_9;
    preRoundConstStage_addContextDelayed_stateElements_10 <= preRoundConstStage_input_payload_delay_16_stateElements_10;
    preRoundConstStage_addContextDelayed_stateElement <= preRoundConstStage_input_payload_delay_16_stateElement;
    if(demuxInst_io_output0_ready) begin
      demuxInst_io_output0_rData_isFull <= demuxInst_io_output0_payload_isFull;
      demuxInst_io_output0_rData_fullRound <= demuxInst_io_output0_payload_fullRound;
      demuxInst_io_output0_rData_partialRound <= demuxInst_io_output0_payload_partialRound;
      demuxInst_io_output0_rData_stateSize <= demuxInst_io_output0_payload_stateSize;
      demuxInst_io_output0_rData_stateID <= demuxInst_io_output0_payload_stateID;
      demuxInst_io_output0_rData_stateElements_0 <= demuxInst_io_output0_payload_stateElements_0;
      demuxInst_io_output0_rData_stateElements_1 <= demuxInst_io_output0_payload_stateElements_1;
      demuxInst_io_output0_rData_stateElements_2 <= demuxInst_io_output0_payload_stateElements_2;
      demuxInst_io_output0_rData_stateElements_3 <= demuxInst_io_output0_payload_stateElements_3;
      demuxInst_io_output0_rData_stateElements_4 <= demuxInst_io_output0_payload_stateElements_4;
      demuxInst_io_output0_rData_stateElements_5 <= demuxInst_io_output0_payload_stateElements_5;
      demuxInst_io_output0_rData_stateElements_6 <= demuxInst_io_output0_payload_stateElements_6;
      demuxInst_io_output0_rData_stateElements_7 <= demuxInst_io_output0_payload_stateElements_7;
      demuxInst_io_output0_rData_stateElements_8 <= demuxInst_io_output0_payload_stateElements_8;
      demuxInst_io_output0_rData_stateElements_9 <= demuxInst_io_output0_payload_stateElements_9;
      demuxInst_io_output0_rData_stateElements_10 <= demuxInst_io_output0_payload_stateElements_10;
      demuxInst_io_output0_rData_stateElements_11 <= demuxInst_io_output0_payload_stateElements_11;
    end
    if(demuxInst_io_output0_s2mPipe_ready) begin
      demuxInst_io_output0_s2mPipe_rData_isFull <= demuxInst_io_output0_s2mPipe_payload_isFull;
      demuxInst_io_output0_s2mPipe_rData_fullRound <= demuxInst_io_output0_s2mPipe_payload_fullRound;
      demuxInst_io_output0_s2mPipe_rData_partialRound <= demuxInst_io_output0_s2mPipe_payload_partialRound;
      demuxInst_io_output0_s2mPipe_rData_stateSize <= demuxInst_io_output0_s2mPipe_payload_stateSize;
      demuxInst_io_output0_s2mPipe_rData_stateID <= demuxInst_io_output0_s2mPipe_payload_stateID;
      demuxInst_io_output0_s2mPipe_rData_stateElements_0 <= demuxInst_io_output0_s2mPipe_payload_stateElements_0;
      demuxInst_io_output0_s2mPipe_rData_stateElements_1 <= demuxInst_io_output0_s2mPipe_payload_stateElements_1;
      demuxInst_io_output0_s2mPipe_rData_stateElements_2 <= demuxInst_io_output0_s2mPipe_payload_stateElements_2;
      demuxInst_io_output0_s2mPipe_rData_stateElements_3 <= demuxInst_io_output0_s2mPipe_payload_stateElements_3;
      demuxInst_io_output0_s2mPipe_rData_stateElements_4 <= demuxInst_io_output0_s2mPipe_payload_stateElements_4;
      demuxInst_io_output0_s2mPipe_rData_stateElements_5 <= demuxInst_io_output0_s2mPipe_payload_stateElements_5;
      demuxInst_io_output0_s2mPipe_rData_stateElements_6 <= demuxInst_io_output0_s2mPipe_payload_stateElements_6;
      demuxInst_io_output0_s2mPipe_rData_stateElements_7 <= demuxInst_io_output0_s2mPipe_payload_stateElements_7;
      demuxInst_io_output0_s2mPipe_rData_stateElements_8 <= demuxInst_io_output0_s2mPipe_payload_stateElements_8;
      demuxInst_io_output0_s2mPipe_rData_stateElements_9 <= demuxInst_io_output0_s2mPipe_payload_stateElements_9;
      demuxInst_io_output0_s2mPipe_rData_stateElements_10 <= demuxInst_io_output0_s2mPipe_payload_stateElements_10;
      demuxInst_io_output0_s2mPipe_rData_stateElements_11 <= demuxInst_io_output0_s2mPipe_payload_stateElements_11;
    end
    if(demuxInst_io_output1_ready) begin
      demuxInst_io_output1_rData_stateID <= demuxInst_io_output1_payload_stateID;
      demuxInst_io_output1_rData_stateElement <= demuxInst_io_output1_payload_stateElement;
    end
  end

  always @(posedge clk) begin
    if(!resetn) begin
      demuxInst_io_output0_rValid <= 1'b0;
      demuxInst_io_output0_s2mPipe_rValid <= 1'b0;
      demuxInst_io_output1_rValid <= 1'b0;
    end else begin
      if(demuxInst_io_output0_valid) begin
        demuxInst_io_output0_rValid <= 1'b1;
      end
      if(demuxInst_io_output0_s2mPipe_ready) begin
        demuxInst_io_output0_rValid <= 1'b0;
      end
      if(demuxInst_io_output0_s2mPipe_ready) begin
        demuxInst_io_output0_s2mPipe_rValid <= demuxInst_io_output0_s2mPipe_valid;
      end
      if(demuxInst_io_output1_ready) begin
        demuxInst_io_output1_rValid <= demuxInst_io_output1_valid;
      end
    end
  end


endmodule

module AXI4StreamReceiver (
  input               io_input_valid,
  output reg          io_input_ready,
  input               io_input_last,
  input      [254:0]  io_input_payload,
  output              io_output_valid,
  input               io_output_ready,
  output              io_output_payload_isFull,
  output     [2:0]    io_output_payload_fullRound,
  output     [5:0]    io_output_payload_partialRound,
  output     [3:0]    io_output_payload_stateSize,
  output     [7:0]    io_output_payload_stateID,
  output     [254:0]  io_output_payload_stateElements_0,
  output     [254:0]  io_output_payload_stateElements_1,
  output     [254:0]  io_output_payload_stateElements_2,
  output     [254:0]  io_output_payload_stateElements_3,
  output     [254:0]  io_output_payload_stateElements_4,
  output     [254:0]  io_output_payload_stateElements_5,
  output     [254:0]  io_output_payload_stateElements_6,
  output     [254:0]  io_output_payload_stateElements_7,
  output     [254:0]  io_output_payload_stateElements_8,
  output     [254:0]  io_output_payload_stateElements_9,
  output     [254:0]  io_output_payload_stateElements_10,
  output     [254:0]  io_output_payload_stateElements_11,
  input               clk,
  input               resetn
);
  localparam receiver_receiverFSM_enumDef_BOOT = 2'd0;
  localparam receiver_receiverFSM_enumDef_BUSY = 2'd1;
  localparam receiver_receiverFSM_enumDef_DONE = 2'd2;

  reg                 receiver_output_valid;
  reg                 receiver_output_ready;
  wire                receiver_output_payload_isFull;
  wire       [2:0]    receiver_output_payload_fullRound;
  wire       [5:0]    receiver_output_payload_partialRound;
  reg        [3:0]    receiver_output_payload_stateSize;
  reg        [7:0]    receiver_output_payload_stateID;
  reg        [254:0]  receiver_output_payload_stateElements_0;
  reg        [254:0]  receiver_output_payload_stateElements_1;
  reg        [254:0]  receiver_output_payload_stateElements_2;
  reg        [254:0]  receiver_output_payload_stateElements_3;
  reg        [254:0]  receiver_output_payload_stateElements_4;
  reg        [254:0]  receiver_output_payload_stateElements_5;
  reg        [254:0]  receiver_output_payload_stateElements_6;
  reg        [254:0]  receiver_output_payload_stateElements_7;
  reg        [254:0]  receiver_output_payload_stateElements_8;
  reg        [254:0]  receiver_output_payload_stateElements_9;
  reg        [254:0]  receiver_output_payload_stateElements_10;
  reg        [254:0]  receiver_output_payload_stateElements_11;
  reg        [3:0]    receiver_sizeCounter;
  reg        [7:0]    receiver_idCounter;
  reg        [254:0]  receiver_buffer_0;
  reg        [254:0]  receiver_buffer_1;
  reg        [254:0]  receiver_buffer_2;
  reg        [254:0]  receiver_buffer_3;
  reg        [254:0]  receiver_buffer_4;
  reg        [254:0]  receiver_buffer_5;
  reg        [254:0]  receiver_buffer_6;
  reg        [254:0]  receiver_buffer_7;
  reg        [254:0]  receiver_buffer_8;
  reg        [254:0]  receiver_buffer_9;
  reg        [254:0]  receiver_buffer_10;
  reg        [254:0]  receiver_buffer_11;
  wire                receiver_receiverFSM_wantExit;
  reg                 receiver_receiverFSM_wantStart;
  wire                receiver_receiverFSM_wantKill;
  wire                receiver_output_m2sPipe_valid;
  wire                receiver_output_m2sPipe_ready;
  wire                receiver_output_m2sPipe_payload_isFull;
  wire       [2:0]    receiver_output_m2sPipe_payload_fullRound;
  wire       [5:0]    receiver_output_m2sPipe_payload_partialRound;
  wire       [3:0]    receiver_output_m2sPipe_payload_stateSize;
  wire       [7:0]    receiver_output_m2sPipe_payload_stateID;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_0;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_1;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_2;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_3;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_4;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_5;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_6;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_7;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_8;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_9;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_10;
  wire       [254:0]  receiver_output_m2sPipe_payload_stateElements_11;
  reg                 receiver_output_rValid;
  reg                 receiver_output_rData_isFull;
  reg        [2:0]    receiver_output_rData_fullRound;
  reg        [5:0]    receiver_output_rData_partialRound;
  reg        [3:0]    receiver_output_rData_stateSize;
  reg        [7:0]    receiver_output_rData_stateID;
  reg        [254:0]  receiver_output_rData_stateElements_0;
  reg        [254:0]  receiver_output_rData_stateElements_1;
  reg        [254:0]  receiver_output_rData_stateElements_2;
  reg        [254:0]  receiver_output_rData_stateElements_3;
  reg        [254:0]  receiver_output_rData_stateElements_4;
  reg        [254:0]  receiver_output_rData_stateElements_5;
  reg        [254:0]  receiver_output_rData_stateElements_6;
  reg        [254:0]  receiver_output_rData_stateElements_7;
  reg        [254:0]  receiver_output_rData_stateElements_8;
  reg        [254:0]  receiver_output_rData_stateElements_9;
  reg        [254:0]  receiver_output_rData_stateElements_10;
  reg        [254:0]  receiver_output_rData_stateElements_11;
  wire                when_Stream_l342;
  reg        [1:0]    receiver_receiverFSM_stateReg;
  reg        [1:0]    receiver_receiverFSM_stateNext;
  wire                when_AXI4StreamInterface_l47;
  wire       [15:0]   _zz_1;
  wire                receiver_output_fire;
  wire                when_AXI4StreamInterface_l67;
  `ifndef SYNTHESIS
  reg [31:0] receiver_receiverFSM_stateReg_string;
  reg [31:0] receiver_receiverFSM_stateNext_string;
  `endif


  `ifndef SYNTHESIS
  always @(*) begin
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BOOT : receiver_receiverFSM_stateReg_string = "BOOT";
      receiver_receiverFSM_enumDef_BUSY : receiver_receiverFSM_stateReg_string = "BUSY";
      receiver_receiverFSM_enumDef_DONE : receiver_receiverFSM_stateReg_string = "DONE";
      default : receiver_receiverFSM_stateReg_string = "????";
    endcase
  end
  always @(*) begin
    case(receiver_receiverFSM_stateNext)
      receiver_receiverFSM_enumDef_BOOT : receiver_receiverFSM_stateNext_string = "BOOT";
      receiver_receiverFSM_enumDef_BUSY : receiver_receiverFSM_stateNext_string = "BUSY";
      receiver_receiverFSM_enumDef_DONE : receiver_receiverFSM_stateNext_string = "DONE";
      default : receiver_receiverFSM_stateNext_string = "????";
    endcase
  end
  `endif

  assign receiver_receiverFSM_wantExit = 1'b0;
  always @(*) begin
    receiver_receiverFSM_wantStart = 1'b0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
      end
      default : begin
        receiver_receiverFSM_wantStart = 1'b1;
      end
    endcase
  end

  assign receiver_receiverFSM_wantKill = 1'b0;
  always @(*) begin
    io_input_ready = 1'b0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
        io_input_ready = 1'b1;
      end
      receiver_receiverFSM_enumDef_DONE : begin
        if(receiver_output_fire) begin
          io_input_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_valid = 1'b0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign receiver_output_payload_isFull = 1'b1;
  assign receiver_output_payload_fullRound = 3'b000;
  assign receiver_output_payload_partialRound = 6'h3f;
  always @(*) begin
    receiver_output_payload_stateSize = 4'b0000;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateSize = receiver_sizeCounter;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateID = 8'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateID = receiver_idCounter;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_0 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_0 = receiver_buffer_0;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_1 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_1 = receiver_buffer_1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_2 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_2 = receiver_buffer_2;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_3 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_3 = receiver_buffer_3;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_4 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_4 = receiver_buffer_4;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_5 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_5 = receiver_buffer_5;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_6 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_6 = receiver_buffer_6;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_7 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_7 = receiver_buffer_7;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_8 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_8 = receiver_buffer_8;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_9 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_9 = receiver_buffer_9;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_10 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_10 = receiver_buffer_10;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_payload_stateElements_11 = 255'h0;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
      end
      receiver_receiverFSM_enumDef_DONE : begin
        receiver_output_payload_stateElements_11 = receiver_buffer_11;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    receiver_output_ready = receiver_output_m2sPipe_ready;
    if(when_Stream_l342) begin
      receiver_output_ready = 1'b1;
    end
  end

  assign when_Stream_l342 = (! receiver_output_m2sPipe_valid);
  assign receiver_output_m2sPipe_valid = receiver_output_rValid;
  assign receiver_output_m2sPipe_payload_isFull = receiver_output_rData_isFull;
  assign receiver_output_m2sPipe_payload_fullRound = receiver_output_rData_fullRound;
  assign receiver_output_m2sPipe_payload_partialRound = receiver_output_rData_partialRound;
  assign receiver_output_m2sPipe_payload_stateSize = receiver_output_rData_stateSize;
  assign receiver_output_m2sPipe_payload_stateID = receiver_output_rData_stateID;
  assign receiver_output_m2sPipe_payload_stateElements_0 = receiver_output_rData_stateElements_0;
  assign receiver_output_m2sPipe_payload_stateElements_1 = receiver_output_rData_stateElements_1;
  assign receiver_output_m2sPipe_payload_stateElements_2 = receiver_output_rData_stateElements_2;
  assign receiver_output_m2sPipe_payload_stateElements_3 = receiver_output_rData_stateElements_3;
  assign receiver_output_m2sPipe_payload_stateElements_4 = receiver_output_rData_stateElements_4;
  assign receiver_output_m2sPipe_payload_stateElements_5 = receiver_output_rData_stateElements_5;
  assign receiver_output_m2sPipe_payload_stateElements_6 = receiver_output_rData_stateElements_6;
  assign receiver_output_m2sPipe_payload_stateElements_7 = receiver_output_rData_stateElements_7;
  assign receiver_output_m2sPipe_payload_stateElements_8 = receiver_output_rData_stateElements_8;
  assign receiver_output_m2sPipe_payload_stateElements_9 = receiver_output_rData_stateElements_9;
  assign receiver_output_m2sPipe_payload_stateElements_10 = receiver_output_rData_stateElements_10;
  assign receiver_output_m2sPipe_payload_stateElements_11 = receiver_output_rData_stateElements_11;
  assign io_output_valid = receiver_output_m2sPipe_valid;
  assign receiver_output_m2sPipe_ready = io_output_ready;
  assign io_output_payload_isFull = receiver_output_m2sPipe_payload_isFull;
  assign io_output_payload_fullRound = receiver_output_m2sPipe_payload_fullRound;
  assign io_output_payload_partialRound = receiver_output_m2sPipe_payload_partialRound;
  assign io_output_payload_stateSize = receiver_output_m2sPipe_payload_stateSize;
  assign io_output_payload_stateID = receiver_output_m2sPipe_payload_stateID;
  assign io_output_payload_stateElements_0 = receiver_output_m2sPipe_payload_stateElements_0;
  assign io_output_payload_stateElements_1 = receiver_output_m2sPipe_payload_stateElements_1;
  assign io_output_payload_stateElements_2 = receiver_output_m2sPipe_payload_stateElements_2;
  assign io_output_payload_stateElements_3 = receiver_output_m2sPipe_payload_stateElements_3;
  assign io_output_payload_stateElements_4 = receiver_output_m2sPipe_payload_stateElements_4;
  assign io_output_payload_stateElements_5 = receiver_output_m2sPipe_payload_stateElements_5;
  assign io_output_payload_stateElements_6 = receiver_output_m2sPipe_payload_stateElements_6;
  assign io_output_payload_stateElements_7 = receiver_output_m2sPipe_payload_stateElements_7;
  assign io_output_payload_stateElements_8 = receiver_output_m2sPipe_payload_stateElements_8;
  assign io_output_payload_stateElements_9 = receiver_output_m2sPipe_payload_stateElements_9;
  assign io_output_payload_stateElements_10 = receiver_output_m2sPipe_payload_stateElements_10;
  assign io_output_payload_stateElements_11 = receiver_output_m2sPipe_payload_stateElements_11;
  always @(*) begin
    receiver_receiverFSM_stateNext = receiver_receiverFSM_stateReg;
    case(receiver_receiverFSM_stateReg)
      receiver_receiverFSM_enumDef_BUSY : begin
        if(when_AXI4StreamInterface_l47) begin
          if(io_input_last) begin
            receiver_receiverFSM_stateNext = receiver_receiverFSM_enumDef_DONE;
          end
        end
      end
      receiver_receiverFSM_enumDef_DONE : begin
        if(receiver_output_fire) begin
          receiver_receiverFSM_stateNext = receiver_receiverFSM_enumDef_BUSY;
        end
      end
      default : begin
      end
    endcase
    if(receiver_receiverFSM_wantStart) begin
      receiver_receiverFSM_stateNext = receiver_receiverFSM_enumDef_BUSY;
    end
    if(receiver_receiverFSM_wantKill) begin
      receiver_receiverFSM_stateNext = receiver_receiverFSM_enumDef_BOOT;
    end
  end

  assign when_AXI4StreamInterface_l47 = (io_input_valid && io_input_ready);
  assign _zz_1 = ({15'd0,1'b1} <<< receiver_sizeCounter);
  assign receiver_output_fire = (receiver_output_valid && receiver_output_ready);
  assign when_AXI4StreamInterface_l67 = (io_input_valid && io_input_ready);
  always @(posedge clk) begin
    if(!resetn) begin
      receiver_sizeCounter <= 4'b0000;
      receiver_idCounter <= 8'h0;
      receiver_buffer_0 <= 255'h0;
      receiver_buffer_1 <= 255'h0;
      receiver_buffer_2 <= 255'h0;
      receiver_buffer_3 <= 255'h0;
      receiver_buffer_4 <= 255'h0;
      receiver_buffer_5 <= 255'h0;
      receiver_buffer_6 <= 255'h0;
      receiver_buffer_7 <= 255'h0;
      receiver_buffer_8 <= 255'h0;
      receiver_buffer_9 <= 255'h0;
      receiver_buffer_10 <= 255'h0;
      receiver_buffer_11 <= 255'h0;
      receiver_output_rValid <= 1'b0;
      receiver_receiverFSM_stateReg <= receiver_receiverFSM_enumDef_BOOT;
    end else begin
      if(receiver_output_ready) begin
        receiver_output_rValid <= receiver_output_valid;
      end
      receiver_receiverFSM_stateReg <= receiver_receiverFSM_stateNext;
      case(receiver_receiverFSM_stateReg)
        receiver_receiverFSM_enumDef_BUSY : begin
          if(when_AXI4StreamInterface_l47) begin
            if(_zz_1[0]) begin
              receiver_buffer_0 <= io_input_payload;
            end
            if(_zz_1[1]) begin
              receiver_buffer_1 <= io_input_payload;
            end
            if(_zz_1[2]) begin
              receiver_buffer_2 <= io_input_payload;
            end
            if(_zz_1[3]) begin
              receiver_buffer_3 <= io_input_payload;
            end
            if(_zz_1[4]) begin
              receiver_buffer_4 <= io_input_payload;
            end
            if(_zz_1[5]) begin
              receiver_buffer_5 <= io_input_payload;
            end
            if(_zz_1[6]) begin
              receiver_buffer_6 <= io_input_payload;
            end
            if(_zz_1[7]) begin
              receiver_buffer_7 <= io_input_payload;
            end
            if(_zz_1[8]) begin
              receiver_buffer_8 <= io_input_payload;
            end
            if(_zz_1[9]) begin
              receiver_buffer_9 <= io_input_payload;
            end
            if(_zz_1[10]) begin
              receiver_buffer_10 <= io_input_payload;
            end
            if(_zz_1[11]) begin
              receiver_buffer_11 <= io_input_payload;
            end
            receiver_sizeCounter <= (receiver_sizeCounter + 4'b0001);
          end
        end
        receiver_receiverFSM_enumDef_DONE : begin
          if(receiver_output_fire) begin
            receiver_buffer_0 <= 255'h0;
            receiver_buffer_1 <= 255'h0;
            receiver_buffer_2 <= 255'h0;
            receiver_buffer_3 <= 255'h0;
            receiver_buffer_4 <= 255'h0;
            receiver_buffer_5 <= 255'h0;
            receiver_buffer_6 <= 255'h0;
            receiver_buffer_7 <= 255'h0;
            receiver_buffer_8 <= 255'h0;
            receiver_buffer_9 <= 255'h0;
            receiver_buffer_10 <= 255'h0;
            receiver_buffer_11 <= 255'h0;
            receiver_idCounter <= (receiver_idCounter + 8'h01);
            receiver_sizeCounter <= 4'b0000;
            if(when_AXI4StreamInterface_l67) begin
              receiver_buffer_0 <= io_input_payload;
              receiver_sizeCounter <= 4'b0001;
            end
          end
        end
        default : begin
        end
      endcase
    end
  end

  always @(posedge clk) begin
    if(receiver_output_ready) begin
      receiver_output_rData_isFull <= receiver_output_payload_isFull;
      receiver_output_rData_fullRound <= receiver_output_payload_fullRound;
      receiver_output_rData_partialRound <= receiver_output_payload_partialRound;
      receiver_output_rData_stateSize <= receiver_output_payload_stateSize;
      receiver_output_rData_stateID <= receiver_output_payload_stateID;
      receiver_output_rData_stateElements_0 <= receiver_output_payload_stateElements_0;
      receiver_output_rData_stateElements_1 <= receiver_output_payload_stateElements_1;
      receiver_output_rData_stateElements_2 <= receiver_output_payload_stateElements_2;
      receiver_output_rData_stateElements_3 <= receiver_output_payload_stateElements_3;
      receiver_output_rData_stateElements_4 <= receiver_output_payload_stateElements_4;
      receiver_output_rData_stateElements_5 <= receiver_output_payload_stateElements_5;
      receiver_output_rData_stateElements_6 <= receiver_output_payload_stateElements_6;
      receiver_output_rData_stateElements_7 <= receiver_output_payload_stateElements_7;
      receiver_output_rData_stateElements_8 <= receiver_output_payload_stateElements_8;
      receiver_output_rData_stateElements_9 <= receiver_output_payload_stateElements_9;
      receiver_output_rData_stateElements_10 <= receiver_output_payload_stateElements_10;
      receiver_output_rData_stateElements_11 <= receiver_output_payload_stateElements_11;
    end
  end


endmodule

module StreamFifo_1 (
  input               io_push_valid,
  output              io_push_ready,
  input      [7:0]    io_push_payload_stateID,
  input      [254:0]  io_push_payload_stateElement,
  output              io_pop_valid,
  input               io_pop_ready,
  output     [7:0]    io_pop_payload_stateID,
  output     [254:0]  io_pop_payload_stateElement,
  input               io_flush,
  output     [3:0]    io_occupancy,
  output     [3:0]    io_availability,
  input               clk,
  input               resetn
);

  reg        [262:0]  _zz_logic_ram_port0;
  wire       [2:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [2:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz__zz_io_pop_payload_stateID;
  wire       [262:0]  _zz_logic_ram_port_1;
  wire       [2:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [2:0]    logic_pushPtr_valueNext;
  reg        [2:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [2:0]    logic_popPtr_valueNext;
  reg        [2:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire       [262:0]  _zz_io_pop_payload_stateID;
  wire                when_Stream_l954;
  wire       [2:0]    logic_ptrDif;
  reg [262:0] logic_ram [0:7];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {2'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {2'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz__zz_io_pop_payload_stateID = 1'b1;
  assign _zz_logic_ram_port_1 = {io_push_payload_stateElement,io_push_payload_stateID};
  always @(posedge clk) begin
    if(_zz__zz_io_pop_payload_stateID) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 3'b111);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 3'b000;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 3'b111);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 3'b000;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign _zz_io_pop_payload_stateID = _zz_logic_ram_port0;
  assign io_pop_payload_stateID = _zz_io_pop_payload_stateID[7 : 0];
  assign io_pop_payload_stateElement = _zz_io_pop_payload_stateID[262 : 8];
  assign when_Stream_l954 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk) begin
    if(!resetn) begin
      logic_pushPtr_value <= 3'b000;
      logic_popPtr_value <= 3'b000;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l954) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module StreamDemux_1 (
  input      [0:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElement,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output     [7:0]    io_outputs_0_payload_stateID,
  output     [254:0]  io_outputs_0_payload_stateElement,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output     [7:0]    io_outputs_1_payload_stateID,
  output     [254:0]  io_outputs_1_payload_stateElement
);

  wire                when_Stream_l764;
  wire                when_Stream_l764_1;

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l764) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l764_1) begin
      io_input_ready = io_outputs_1_ready;
    end
  end

  assign io_outputs_0_payload_stateID = io_input_payload_stateID;
  assign io_outputs_0_payload_stateElement = io_input_payload_stateElement;
  assign when_Stream_l764 = (1'b0 != io_select);
  always @(*) begin
    if(when_Stream_l764) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_stateID = io_input_payload_stateID;
  assign io_outputs_1_payload_stateElement = io_input_payload_stateElement;
  assign when_Stream_l764_1 = (1'b1 != io_select);
  always @(*) begin
    if(when_Stream_l764_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end


endmodule

module StreamArbiter_1 (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input      [7:0]    io_inputs_0_payload_stateID,
  input      [254:0]  io_inputs_0_payload_stateElement,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input      [7:0]    io_inputs_1_payload_stateID,
  input      [254:0]  io_inputs_1_payload_stateElement,
  output              io_output_valid,
  input               io_output_ready,
  output     [7:0]    io_output_payload_stateID,
  output     [254:0]  io_output_payload_stateElement,
  output     [0:0]    io_chosen,
  output     [1:0]    io_chosenOH,
  input               clk,
  input               resetn
);

  wire       [1:0]    _zz_maskProposal_1_1;
  wire       [1:0]    _zz_maskProposal_1_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_1;
  wire                io_output_fire;
  wire                _zz_io_chosen;

  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz_maskProposal_1_2));
  assign _zz_maskProposal_1_2 = (_zz_maskProposal_1 - 2'b01);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_1 = {io_inputs_1_valid,io_inputs_0_valid};
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_stateID = (maskRouted_0 ? io_inputs_0_payload_stateID : io_inputs_1_payload_stateID);
  assign io_output_payload_stateElement = (maskRouted_0 ? io_inputs_0_payload_stateElement : io_inputs_1_payload_stateElement);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk) begin
    if(!resetn) begin
      locked <= 1'b0;
    end else begin
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
    end
  end


endmodule

module BundleFifo (
  input               io_push_valid,
  output              io_push_ready,
  input               io_push_payload_isFull,
  input      [2:0]    io_push_payload_fullRound,
  input      [5:0]    io_push_payload_partialRound,
  input      [3:0]    io_push_payload_stateSize,
  input      [7:0]    io_push_payload_stateID,
  input      [254:0]  io_push_payload_stateElements_0,
  input      [254:0]  io_push_payload_stateElements_1,
  input      [254:0]  io_push_payload_stateElements_2,
  input      [254:0]  io_push_payload_stateElements_3,
  input      [254:0]  io_push_payload_stateElements_4,
  input      [254:0]  io_push_payload_stateElements_5,
  input      [254:0]  io_push_payload_stateElements_6,
  input      [254:0]  io_push_payload_stateElements_7,
  input      [254:0]  io_push_payload_stateElements_8,
  input      [254:0]  io_push_payload_stateElements_9,
  input      [254:0]  io_push_payload_stateElements_10,
  input      [254:0]  io_push_payload_stateElements_11,
  output              io_pop_valid,
  input               io_pop_ready,
  output              io_pop_payload_isFull,
  output     [2:0]    io_pop_payload_fullRound,
  output     [5:0]    io_pop_payload_partialRound,
  output     [3:0]    io_pop_payload_stateSize,
  output     [7:0]    io_pop_payload_stateID,
  output     [254:0]  io_pop_payload_stateElements_0,
  output     [254:0]  io_pop_payload_stateElements_1,
  output     [254:0]  io_pop_payload_stateElements_2,
  output     [254:0]  io_pop_payload_stateElements_3,
  output     [254:0]  io_pop_payload_stateElements_4,
  output     [254:0]  io_pop_payload_stateElements_5,
  output     [254:0]  io_pop_payload_stateElements_6,
  output     [254:0]  io_pop_payload_stateElements_7,
  output     [254:0]  io_pop_payload_stateElements_8,
  output     [254:0]  io_pop_payload_stateElements_9,
  output     [254:0]  io_pop_payload_stateElements_10,
  output     [254:0]  io_pop_payload_stateElements_11,
  input               clk,
  input               resetn
);

  wire                io_push_fifo_io_push_ready;
  wire                io_push_fifo_io_pop_valid;
  wire                io_push_fifo_io_pop_payload_isFull;
  wire       [2:0]    io_push_fifo_io_pop_payload_fullRound;
  wire       [5:0]    io_push_fifo_io_pop_payload_partialRound;
  wire       [3:0]    io_push_fifo_io_pop_payload_stateSize;
  wire       [7:0]    io_push_fifo_io_pop_payload_stateID;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_0;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_1;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_2;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_3;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_4;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_5;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_6;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_7;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_8;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_9;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_10;
  wire       [254:0]  io_push_fifo_io_pop_payload_stateElements_11;
  wire       [8:0]    io_push_fifo_io_occupancy;
  wire       [8:0]    io_push_fifo_io_availability;

  StreamFifo io_push_fifo (
    .io_push_valid                       (io_push_valid                                        ), //i
    .io_push_ready                       (io_push_fifo_io_push_ready                           ), //o
    .io_push_payload_isFull              (io_push_payload_isFull                               ), //i
    .io_push_payload_fullRound           (io_push_payload_fullRound[2:0]                       ), //i
    .io_push_payload_partialRound        (io_push_payload_partialRound[5:0]                    ), //i
    .io_push_payload_stateSize           (io_push_payload_stateSize[3:0]                       ), //i
    .io_push_payload_stateID             (io_push_payload_stateID[7:0]                         ), //i
    .io_push_payload_stateElements_0     (io_push_payload_stateElements_0[254:0]               ), //i
    .io_push_payload_stateElements_1     (io_push_payload_stateElements_1[254:0]               ), //i
    .io_push_payload_stateElements_2     (io_push_payload_stateElements_2[254:0]               ), //i
    .io_push_payload_stateElements_3     (io_push_payload_stateElements_3[254:0]               ), //i
    .io_push_payload_stateElements_4     (io_push_payload_stateElements_4[254:0]               ), //i
    .io_push_payload_stateElements_5     (io_push_payload_stateElements_5[254:0]               ), //i
    .io_push_payload_stateElements_6     (io_push_payload_stateElements_6[254:0]               ), //i
    .io_push_payload_stateElements_7     (io_push_payload_stateElements_7[254:0]               ), //i
    .io_push_payload_stateElements_8     (io_push_payload_stateElements_8[254:0]               ), //i
    .io_push_payload_stateElements_9     (io_push_payload_stateElements_9[254:0]               ), //i
    .io_push_payload_stateElements_10    (io_push_payload_stateElements_10[254:0]              ), //i
    .io_push_payload_stateElements_11    (io_push_payload_stateElements_11[254:0]              ), //i
    .io_pop_valid                        (io_push_fifo_io_pop_valid                            ), //o
    .io_pop_ready                        (io_pop_ready                                         ), //i
    .io_pop_payload_isFull               (io_push_fifo_io_pop_payload_isFull                   ), //o
    .io_pop_payload_fullRound            (io_push_fifo_io_pop_payload_fullRound[2:0]           ), //o
    .io_pop_payload_partialRound         (io_push_fifo_io_pop_payload_partialRound[5:0]        ), //o
    .io_pop_payload_stateSize            (io_push_fifo_io_pop_payload_stateSize[3:0]           ), //o
    .io_pop_payload_stateID              (io_push_fifo_io_pop_payload_stateID[7:0]             ), //o
    .io_pop_payload_stateElements_0      (io_push_fifo_io_pop_payload_stateElements_0[254:0]   ), //o
    .io_pop_payload_stateElements_1      (io_push_fifo_io_pop_payload_stateElements_1[254:0]   ), //o
    .io_pop_payload_stateElements_2      (io_push_fifo_io_pop_payload_stateElements_2[254:0]   ), //o
    .io_pop_payload_stateElements_3      (io_push_fifo_io_pop_payload_stateElements_3[254:0]   ), //o
    .io_pop_payload_stateElements_4      (io_push_fifo_io_pop_payload_stateElements_4[254:0]   ), //o
    .io_pop_payload_stateElements_5      (io_push_fifo_io_pop_payload_stateElements_5[254:0]   ), //o
    .io_pop_payload_stateElements_6      (io_push_fifo_io_pop_payload_stateElements_6[254:0]   ), //o
    .io_pop_payload_stateElements_7      (io_push_fifo_io_pop_payload_stateElements_7[254:0]   ), //o
    .io_pop_payload_stateElements_8      (io_push_fifo_io_pop_payload_stateElements_8[254:0]   ), //o
    .io_pop_payload_stateElements_9      (io_push_fifo_io_pop_payload_stateElements_9[254:0]   ), //o
    .io_pop_payload_stateElements_10     (io_push_fifo_io_pop_payload_stateElements_10[254:0]  ), //o
    .io_pop_payload_stateElements_11     (io_push_fifo_io_pop_payload_stateElements_11[254:0]  ), //o
    .io_flush                            (1'b0                                                 ), //i
    .io_occupancy                        (io_push_fifo_io_occupancy[8:0]                       ), //o
    .io_availability                     (io_push_fifo_io_availability[8:0]                    ), //o
    .clk                                 (clk                                                  ), //i
    .resetn                              (resetn                                               )  //i
  );
  assign io_push_ready = io_push_fifo_io_push_ready;
  assign io_pop_valid = io_push_fifo_io_pop_valid;
  assign io_pop_payload_isFull = io_push_fifo_io_pop_payload_isFull;
  assign io_pop_payload_fullRound = io_push_fifo_io_pop_payload_fullRound;
  assign io_pop_payload_partialRound = io_push_fifo_io_pop_payload_partialRound;
  assign io_pop_payload_stateSize = io_push_fifo_io_pop_payload_stateSize;
  assign io_pop_payload_stateID = io_push_fifo_io_pop_payload_stateID;
  assign io_pop_payload_stateElements_0 = io_push_fifo_io_pop_payload_stateElements_0;
  assign io_pop_payload_stateElements_1 = io_push_fifo_io_pop_payload_stateElements_1;
  assign io_pop_payload_stateElements_2 = io_push_fifo_io_pop_payload_stateElements_2;
  assign io_pop_payload_stateElements_3 = io_push_fifo_io_pop_payload_stateElements_3;
  assign io_pop_payload_stateElements_4 = io_push_fifo_io_pop_payload_stateElements_4;
  assign io_pop_payload_stateElements_5 = io_push_fifo_io_pop_payload_stateElements_5;
  assign io_pop_payload_stateElements_6 = io_push_fifo_io_pop_payload_stateElements_6;
  assign io_pop_payload_stateElements_7 = io_push_fifo_io_pop_payload_stateElements_7;
  assign io_pop_payload_stateElements_8 = io_push_fifo_io_pop_payload_stateElements_8;
  assign io_pop_payload_stateElements_9 = io_push_fifo_io_pop_payload_stateElements_9;
  assign io_pop_payload_stateElements_10 = io_push_fifo_io_pop_payload_stateElements_10;
  assign io_pop_payload_stateElements_11 = io_push_fifo_io_pop_payload_stateElements_11;

endmodule

module LoopbackDeMux (
  input               io_input_valid,
  output              io_input_ready,
  input               io_input_payload_isFull,
  input      [2:0]    io_input_payload_fullRound,
  input      [5:0]    io_input_payload_partialRound,
  input      [3:0]    io_input_payload_stateSize,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElements_0,
  input      [254:0]  io_input_payload_stateElements_1,
  input      [254:0]  io_input_payload_stateElements_2,
  input      [254:0]  io_input_payload_stateElements_3,
  input      [254:0]  io_input_payload_stateElements_4,
  input      [254:0]  io_input_payload_stateElements_5,
  input      [254:0]  io_input_payload_stateElements_6,
  input      [254:0]  io_input_payload_stateElements_7,
  input      [254:0]  io_input_payload_stateElements_8,
  input      [254:0]  io_input_payload_stateElements_9,
  input      [254:0]  io_input_payload_stateElements_10,
  input      [254:0]  io_input_payload_stateElements_11,
  output              io_output0_valid,
  input               io_output0_ready,
  output              io_output0_payload_isFull,
  output     [2:0]    io_output0_payload_fullRound,
  output     [5:0]    io_output0_payload_partialRound,
  output     [3:0]    io_output0_payload_stateSize,
  output     [7:0]    io_output0_payload_stateID,
  output     [254:0]  io_output0_payload_stateElements_0,
  output     [254:0]  io_output0_payload_stateElements_1,
  output     [254:0]  io_output0_payload_stateElements_2,
  output     [254:0]  io_output0_payload_stateElements_3,
  output     [254:0]  io_output0_payload_stateElements_4,
  output     [254:0]  io_output0_payload_stateElements_5,
  output     [254:0]  io_output0_payload_stateElements_6,
  output     [254:0]  io_output0_payload_stateElements_7,
  output     [254:0]  io_output0_payload_stateElements_8,
  output     [254:0]  io_output0_payload_stateElements_9,
  output     [254:0]  io_output0_payload_stateElements_10,
  output     [254:0]  io_output0_payload_stateElements_11,
  output              io_output1_valid,
  input               io_output1_ready,
  output     [7:0]    io_output1_payload_stateID,
  output     [254:0]  io_output1_payload_stateElement
);

  wire       [0:0]    streamDemux_2_io_select;
  wire                streamDemux_2_io_input_ready;
  wire                streamDemux_2_io_outputs_0_valid;
  wire                streamDemux_2_io_outputs_0_payload_isFull;
  wire       [2:0]    streamDemux_2_io_outputs_0_payload_fullRound;
  wire       [5:0]    streamDemux_2_io_outputs_0_payload_partialRound;
  wire       [3:0]    streamDemux_2_io_outputs_0_payload_stateSize;
  wire       [7:0]    streamDemux_2_io_outputs_0_payload_stateID;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_0;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_1;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_2;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_3;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_4;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_5;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_6;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_7;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_8;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_9;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_10;
  wire       [254:0]  streamDemux_2_io_outputs_0_payload_stateElements_11;
  wire                streamDemux_2_io_outputs_1_valid;
  wire                streamDemux_2_io_outputs_1_payload_isFull;
  wire       [2:0]    streamDemux_2_io_outputs_1_payload_fullRound;
  wire       [5:0]    streamDemux_2_io_outputs_1_payload_partialRound;
  wire       [3:0]    streamDemux_2_io_outputs_1_payload_stateSize;
  wire       [7:0]    streamDemux_2_io_outputs_1_payload_stateID;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_0;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_1;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_2;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_3;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_4;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_5;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_6;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_7;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_8;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_9;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_10;
  wire       [254:0]  streamDemux_2_io_outputs_1_payload_stateElements_11;
  wire       [3:0]    _zz__zz_isFull;
  wire       [5:0]    _zz__zz_isFull_1;
  wire                _zz__zz_isFull_2;
  wire                _zz__zz_isFull_3;
  wire                _zz__zz_isFull_4;
  wire                _zz__zz_isFull_5;
  wire       [2:0]    _zz__zz_fullRound;
  wire       [0:0]    _zz__zz_fullRound_1;
  wire       [5:0]    _zz__zz_partialRound;
  wire       [0:0]    _zz__zz_partialRound_1;
  wire                select_1;
  reg                 _zz_isFull;
  reg        [2:0]    _zz_fullRound;
  reg        [5:0]    _zz_partialRound;
  wire                streamDemux_2_io_outputs_0_translated_valid;
  wire                streamDemux_2_io_outputs_0_translated_ready;
  wire                streamDemux_2_io_outputs_0_translated_payload_isFull;
  wire       [2:0]    streamDemux_2_io_outputs_0_translated_payload_fullRound;
  wire       [5:0]    streamDemux_2_io_outputs_0_translated_payload_partialRound;
  wire       [3:0]    streamDemux_2_io_outputs_0_translated_payload_stateSize;
  wire       [7:0]    streamDemux_2_io_outputs_0_translated_payload_stateID;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_0;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_1;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_2;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_3;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_4;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_5;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_6;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_7;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_8;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_9;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_10;
  wire       [254:0]  streamDemux_2_io_outputs_0_translated_payload_stateElements_11;
  wire                streamDemux_2_io_outputs_1_translated_valid;
  wire                streamDemux_2_io_outputs_1_translated_ready;
  wire       [7:0]    streamDemux_2_io_outputs_1_translated_payload_stateID;
  wire       [254:0]  streamDemux_2_io_outputs_1_translated_payload_stateElement;

  assign _zz__zz_fullRound_1 = _zz_isFull;
  assign _zz__zz_fullRound = {2'd0, _zz__zz_fullRound_1};
  assign _zz__zz_partialRound_1 = (! _zz_isFull);
  assign _zz__zz_partialRound = {5'd0, _zz__zz_partialRound_1};
  assign _zz__zz_isFull = 4'b1001;
  assign _zz__zz_isFull_1 = 6'h38;
  assign _zz__zz_isFull_2 = (io_input_payload_stateSize == 4'b0101);
  assign _zz__zz_isFull_3 = (io_input_payload_partialRound == 6'h37);
  assign _zz__zz_isFull_4 = (io_input_payload_stateSize == 4'b0011);
  assign _zz__zz_isFull_5 = (io_input_payload_partialRound == 6'h36);
  StreamDemux streamDemux_2 (
    .io_select                                (streamDemux_2_io_select                                     ), //i
    .io_input_valid                           (io_input_valid                                              ), //i
    .io_input_ready                           (streamDemux_2_io_input_ready                                ), //o
    .io_input_payload_isFull                  (io_input_payload_isFull                                     ), //i
    .io_input_payload_fullRound               (io_input_payload_fullRound[2:0]                             ), //i
    .io_input_payload_partialRound            (io_input_payload_partialRound[5:0]                          ), //i
    .io_input_payload_stateSize               (io_input_payload_stateSize[3:0]                             ), //i
    .io_input_payload_stateID                 (io_input_payload_stateID[7:0]                               ), //i
    .io_input_payload_stateElements_0         (io_input_payload_stateElements_0[254:0]                     ), //i
    .io_input_payload_stateElements_1         (io_input_payload_stateElements_1[254:0]                     ), //i
    .io_input_payload_stateElements_2         (io_input_payload_stateElements_2[254:0]                     ), //i
    .io_input_payload_stateElements_3         (io_input_payload_stateElements_3[254:0]                     ), //i
    .io_input_payload_stateElements_4         (io_input_payload_stateElements_4[254:0]                     ), //i
    .io_input_payload_stateElements_5         (io_input_payload_stateElements_5[254:0]                     ), //i
    .io_input_payload_stateElements_6         (io_input_payload_stateElements_6[254:0]                     ), //i
    .io_input_payload_stateElements_7         (io_input_payload_stateElements_7[254:0]                     ), //i
    .io_input_payload_stateElements_8         (io_input_payload_stateElements_8[254:0]                     ), //i
    .io_input_payload_stateElements_9         (io_input_payload_stateElements_9[254:0]                     ), //i
    .io_input_payload_stateElements_10        (io_input_payload_stateElements_10[254:0]                    ), //i
    .io_input_payload_stateElements_11        (io_input_payload_stateElements_11[254:0]                    ), //i
    .io_outputs_0_valid                       (streamDemux_2_io_outputs_0_valid                            ), //o
    .io_outputs_0_ready                       (streamDemux_2_io_outputs_0_translated_ready                 ), //i
    .io_outputs_0_payload_isFull              (streamDemux_2_io_outputs_0_payload_isFull                   ), //o
    .io_outputs_0_payload_fullRound           (streamDemux_2_io_outputs_0_payload_fullRound[2:0]           ), //o
    .io_outputs_0_payload_partialRound        (streamDemux_2_io_outputs_0_payload_partialRound[5:0]        ), //o
    .io_outputs_0_payload_stateSize           (streamDemux_2_io_outputs_0_payload_stateSize[3:0]           ), //o
    .io_outputs_0_payload_stateID             (streamDemux_2_io_outputs_0_payload_stateID[7:0]             ), //o
    .io_outputs_0_payload_stateElements_0     (streamDemux_2_io_outputs_0_payload_stateElements_0[254:0]   ), //o
    .io_outputs_0_payload_stateElements_1     (streamDemux_2_io_outputs_0_payload_stateElements_1[254:0]   ), //o
    .io_outputs_0_payload_stateElements_2     (streamDemux_2_io_outputs_0_payload_stateElements_2[254:0]   ), //o
    .io_outputs_0_payload_stateElements_3     (streamDemux_2_io_outputs_0_payload_stateElements_3[254:0]   ), //o
    .io_outputs_0_payload_stateElements_4     (streamDemux_2_io_outputs_0_payload_stateElements_4[254:0]   ), //o
    .io_outputs_0_payload_stateElements_5     (streamDemux_2_io_outputs_0_payload_stateElements_5[254:0]   ), //o
    .io_outputs_0_payload_stateElements_6     (streamDemux_2_io_outputs_0_payload_stateElements_6[254:0]   ), //o
    .io_outputs_0_payload_stateElements_7     (streamDemux_2_io_outputs_0_payload_stateElements_7[254:0]   ), //o
    .io_outputs_0_payload_stateElements_8     (streamDemux_2_io_outputs_0_payload_stateElements_8[254:0]   ), //o
    .io_outputs_0_payload_stateElements_9     (streamDemux_2_io_outputs_0_payload_stateElements_9[254:0]   ), //o
    .io_outputs_0_payload_stateElements_10    (streamDemux_2_io_outputs_0_payload_stateElements_10[254:0]  ), //o
    .io_outputs_0_payload_stateElements_11    (streamDemux_2_io_outputs_0_payload_stateElements_11[254:0]  ), //o
    .io_outputs_1_valid                       (streamDemux_2_io_outputs_1_valid                            ), //o
    .io_outputs_1_ready                       (streamDemux_2_io_outputs_1_translated_ready                 ), //i
    .io_outputs_1_payload_isFull              (streamDemux_2_io_outputs_1_payload_isFull                   ), //o
    .io_outputs_1_payload_fullRound           (streamDemux_2_io_outputs_1_payload_fullRound[2:0]           ), //o
    .io_outputs_1_payload_partialRound        (streamDemux_2_io_outputs_1_payload_partialRound[5:0]        ), //o
    .io_outputs_1_payload_stateSize           (streamDemux_2_io_outputs_1_payload_stateSize[3:0]           ), //o
    .io_outputs_1_payload_stateID             (streamDemux_2_io_outputs_1_payload_stateID[7:0]             ), //o
    .io_outputs_1_payload_stateElements_0     (streamDemux_2_io_outputs_1_payload_stateElements_0[254:0]   ), //o
    .io_outputs_1_payload_stateElements_1     (streamDemux_2_io_outputs_1_payload_stateElements_1[254:0]   ), //o
    .io_outputs_1_payload_stateElements_2     (streamDemux_2_io_outputs_1_payload_stateElements_2[254:0]   ), //o
    .io_outputs_1_payload_stateElements_3     (streamDemux_2_io_outputs_1_payload_stateElements_3[254:0]   ), //o
    .io_outputs_1_payload_stateElements_4     (streamDemux_2_io_outputs_1_payload_stateElements_4[254:0]   ), //o
    .io_outputs_1_payload_stateElements_5     (streamDemux_2_io_outputs_1_payload_stateElements_5[254:0]   ), //o
    .io_outputs_1_payload_stateElements_6     (streamDemux_2_io_outputs_1_payload_stateElements_6[254:0]   ), //o
    .io_outputs_1_payload_stateElements_7     (streamDemux_2_io_outputs_1_payload_stateElements_7[254:0]   ), //o
    .io_outputs_1_payload_stateElements_8     (streamDemux_2_io_outputs_1_payload_stateElements_8[254:0]   ), //o
    .io_outputs_1_payload_stateElements_9     (streamDemux_2_io_outputs_1_payload_stateElements_9[254:0]   ), //o
    .io_outputs_1_payload_stateElements_10    (streamDemux_2_io_outputs_1_payload_stateElements_10[254:0]  ), //o
    .io_outputs_1_payload_stateElements_11    (streamDemux_2_io_outputs_1_payload_stateElements_11[254:0]  )  //o
  );
  assign select_1 = (io_input_payload_fullRound == 3'b111);
  assign io_input_ready = streamDemux_2_io_input_ready;
  assign streamDemux_2_io_select = select_1;
  always @(*) begin
    _zz_isFull = io_input_payload_isFull;
    _zz_isFull = ((io_input_payload_fullRound < 3'b011) || (|{((io_input_payload_stateSize == 4'b1100) && (io_input_payload_partialRound == 6'h38)),{((io_input_payload_stateSize == _zz__zz_isFull) && (io_input_payload_partialRound == _zz__zz_isFull_1)),{(_zz__zz_isFull_2 && _zz__zz_isFull_3),(_zz__zz_isFull_4 && _zz__zz_isFull_5)}}}));
  end

  always @(*) begin
    _zz_fullRound = io_input_payload_fullRound;
    _zz_fullRound = (io_input_payload_fullRound + _zz__zz_fullRound);
  end

  always @(*) begin
    _zz_partialRound = io_input_payload_partialRound;
    _zz_partialRound = (io_input_payload_partialRound + _zz__zz_partialRound);
  end

  assign streamDemux_2_io_outputs_0_translated_valid = streamDemux_2_io_outputs_0_valid;
  assign streamDemux_2_io_outputs_0_translated_payload_isFull = _zz_isFull;
  assign streamDemux_2_io_outputs_0_translated_payload_fullRound = _zz_fullRound;
  assign streamDemux_2_io_outputs_0_translated_payload_partialRound = _zz_partialRound;
  assign streamDemux_2_io_outputs_0_translated_payload_stateSize = io_input_payload_stateSize;
  assign streamDemux_2_io_outputs_0_translated_payload_stateID = io_input_payload_stateID;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_0 = io_input_payload_stateElements_0;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_1 = io_input_payload_stateElements_1;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_2 = io_input_payload_stateElements_2;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_3 = io_input_payload_stateElements_3;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_4 = io_input_payload_stateElements_4;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_5 = io_input_payload_stateElements_5;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_6 = io_input_payload_stateElements_6;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_7 = io_input_payload_stateElements_7;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_8 = io_input_payload_stateElements_8;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_9 = io_input_payload_stateElements_9;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_10 = io_input_payload_stateElements_10;
  assign streamDemux_2_io_outputs_0_translated_payload_stateElements_11 = io_input_payload_stateElements_11;
  assign io_output0_valid = streamDemux_2_io_outputs_0_translated_valid;
  assign streamDemux_2_io_outputs_0_translated_ready = io_output0_ready;
  assign io_output0_payload_isFull = streamDemux_2_io_outputs_0_translated_payload_isFull;
  assign io_output0_payload_fullRound = streamDemux_2_io_outputs_0_translated_payload_fullRound;
  assign io_output0_payload_partialRound = streamDemux_2_io_outputs_0_translated_payload_partialRound;
  assign io_output0_payload_stateSize = streamDemux_2_io_outputs_0_translated_payload_stateSize;
  assign io_output0_payload_stateID = streamDemux_2_io_outputs_0_translated_payload_stateID;
  assign io_output0_payload_stateElements_0 = streamDemux_2_io_outputs_0_translated_payload_stateElements_0;
  assign io_output0_payload_stateElements_1 = streamDemux_2_io_outputs_0_translated_payload_stateElements_1;
  assign io_output0_payload_stateElements_2 = streamDemux_2_io_outputs_0_translated_payload_stateElements_2;
  assign io_output0_payload_stateElements_3 = streamDemux_2_io_outputs_0_translated_payload_stateElements_3;
  assign io_output0_payload_stateElements_4 = streamDemux_2_io_outputs_0_translated_payload_stateElements_4;
  assign io_output0_payload_stateElements_5 = streamDemux_2_io_outputs_0_translated_payload_stateElements_5;
  assign io_output0_payload_stateElements_6 = streamDemux_2_io_outputs_0_translated_payload_stateElements_6;
  assign io_output0_payload_stateElements_7 = streamDemux_2_io_outputs_0_translated_payload_stateElements_7;
  assign io_output0_payload_stateElements_8 = streamDemux_2_io_outputs_0_translated_payload_stateElements_8;
  assign io_output0_payload_stateElements_9 = streamDemux_2_io_outputs_0_translated_payload_stateElements_9;
  assign io_output0_payload_stateElements_10 = streamDemux_2_io_outputs_0_translated_payload_stateElements_10;
  assign io_output0_payload_stateElements_11 = streamDemux_2_io_outputs_0_translated_payload_stateElements_11;
  assign streamDemux_2_io_outputs_1_translated_valid = streamDemux_2_io_outputs_1_valid;
  assign streamDemux_2_io_outputs_1_translated_payload_stateID = streamDemux_2_io_outputs_1_payload_stateID;
  assign streamDemux_2_io_outputs_1_translated_payload_stateElement = streamDemux_2_io_outputs_1_payload_stateElements_1;
  assign io_output1_valid = streamDemux_2_io_outputs_1_translated_valid;
  assign streamDemux_2_io_outputs_1_translated_ready = io_output1_ready;
  assign io_output1_payload_stateID = streamDemux_2_io_outputs_1_translated_payload_stateID;
  assign io_output1_payload_stateElement = streamDemux_2_io_outputs_1_translated_payload_stateElement;

endmodule

module PoseidonThread (
  input               io_input_valid,
  input               io_input_payload_isFull,
  input      [2:0]    io_input_payload_fullRound,
  input      [5:0]    io_input_payload_partialRound,
  input      [3:0]    io_input_payload_stateIndex,
  input      [3:0]    io_input_payload_stateSize,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElements_0,
  input      [254:0]  io_input_payload_stateElements_1,
  input      [254:0]  io_input_payload_stateElements_2,
  input      [254:0]  io_input_payload_stateElements_3,
  input      [254:0]  io_input_payload_stateElements_4,
  input      [254:0]  io_input_payload_stateElements_5,
  input      [254:0]  io_input_payload_stateElements_6,
  input      [254:0]  io_input_payload_stateElements_7,
  input      [254:0]  io_input_payload_stateElements_8,
  input      [254:0]  io_input_payload_stateElements_9,
  input      [254:0]  io_input_payload_stateElements_10,
  input      [254:0]  io_input_payload_stateElement,
  output              io_output_valid,
  output              io_output_payload_isFull,
  output     [2:0]    io_output_payload_fullRound,
  output     [5:0]    io_output_payload_partialRound,
  output     [3:0]    io_output_payload_stateSize,
  output     [7:0]    io_output_payload_stateID,
  output     [254:0]  io_output_payload_stateElements_0,
  output     [254:0]  io_output_payload_stateElements_1,
  output     [254:0]  io_output_payload_stateElements_2,
  output     [254:0]  io_output_payload_stateElements_3,
  output     [254:0]  io_output_payload_stateElements_4,
  output     [254:0]  io_output_payload_stateElements_5,
  output     [254:0]  io_output_payload_stateElements_6,
  output     [254:0]  io_output_payload_stateElements_7,
  output     [254:0]  io_output_payload_stateElements_8,
  output     [254:0]  io_output_payload_stateElements_9,
  output     [254:0]  io_output_payload_stateElements_10,
  output     [254:0]  io_output_payload_stateElements_11,
  input               clk,
  input               resetn
);

  wire                SBox5Stage_montMultiplier0_io_output_valid;
  wire       [254:0]  SBox5Stage_montMultiplier0_io_output_payload_res;
  wire                SBox5Stage_montMultiplier1_io_output_valid;
  wire       [254:0]  SBox5Stage_montMultiplier1_io_output_payload_res;
  wire                SBox5Stage_montMultiplier2_io_output_valid;
  wire       [254:0]  SBox5Stage_montMultiplier2_io_output_payload_res;
  wire       [254:0]  AddRoundConstantStage_constantMemory_io_data;
  wire                AddRoundConstantStage_modAdder_io_output_valid;
  wire       [254:0]  AddRoundConstantStage_modAdder_io_output_payload_res;
  wire                mDSMatrixMultiplier_1_io_output_valid;
  wire                mDSMatrixMultiplier_1_io_output_payload_isFull;
  wire       [2:0]    mDSMatrixMultiplier_1_io_output_payload_fullRound;
  wire       [5:0]    mDSMatrixMultiplier_1_io_output_payload_partialRound;
  wire       [3:0]    mDSMatrixMultiplier_1_io_output_payload_stateSize;
  wire       [7:0]    mDSMatrixMultiplier_1_io_output_payload_stateID;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_0;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_1;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_2;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_3;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_4;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_5;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_6;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_7;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_8;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_9;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_10;
  wire       [254:0]  mDSMatrixMultiplier_1_io_output_payload_stateElements_11;
  wire                mDSMatrixAdders_1_io_output_valid;
  wire                mDSMatrixAdders_1_io_output_payload_isFull;
  wire       [2:0]    mDSMatrixAdders_1_io_output_payload_fullRound;
  wire       [5:0]    mDSMatrixAdders_1_io_output_payload_partialRound;
  wire       [3:0]    mDSMatrixAdders_1_io_output_payload_stateSize;
  wire       [7:0]    mDSMatrixAdders_1_io_output_payload_stateID;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_0;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_1;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_2;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_3;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_4;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_5;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_6;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_7;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_8;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_9;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_10;
  wire       [254:0]  mDSMatrixAdders_1_io_output_payload_stateElements_11;
  wire                SBox5Stage_mulInput0_valid;
  wire       [254:0]  SBox5Stage_mulInput0_payload_op1;
  wire       [254:0]  SBox5Stage_mulInput0_payload_op2;
  wire                SBox5Stage_mulInput1_valid;
  wire       [254:0]  SBox5Stage_mulInput1_payload_op1;
  wire       [254:0]  SBox5Stage_mulInput1_payload_op2;
  reg                 io_input_payload_delay_1_isFull;
  reg        [2:0]    io_input_payload_delay_1_fullRound;
  reg        [5:0]    io_input_payload_delay_1_partialRound;
  reg        [3:0]    io_input_payload_delay_1_stateIndex;
  reg        [3:0]    io_input_payload_delay_1_stateSize;
  reg        [7:0]    io_input_payload_delay_1_stateID;
  reg        [254:0]  io_input_payload_delay_1_stateElements_0;
  reg        [254:0]  io_input_payload_delay_1_stateElements_1;
  reg        [254:0]  io_input_payload_delay_1_stateElements_2;
  reg        [254:0]  io_input_payload_delay_1_stateElements_3;
  reg        [254:0]  io_input_payload_delay_1_stateElements_4;
  reg        [254:0]  io_input_payload_delay_1_stateElements_5;
  reg        [254:0]  io_input_payload_delay_1_stateElements_6;
  reg        [254:0]  io_input_payload_delay_1_stateElements_7;
  reg        [254:0]  io_input_payload_delay_1_stateElements_8;
  reg        [254:0]  io_input_payload_delay_1_stateElements_9;
  reg        [254:0]  io_input_payload_delay_1_stateElements_10;
  reg        [254:0]  io_input_payload_delay_1_stateElement;
  reg                 io_input_payload_delay_2_isFull;
  reg        [2:0]    io_input_payload_delay_2_fullRound;
  reg        [5:0]    io_input_payload_delay_2_partialRound;
  reg        [3:0]    io_input_payload_delay_2_stateIndex;
  reg        [3:0]    io_input_payload_delay_2_stateSize;
  reg        [7:0]    io_input_payload_delay_2_stateID;
  reg        [254:0]  io_input_payload_delay_2_stateElements_0;
  reg        [254:0]  io_input_payload_delay_2_stateElements_1;
  reg        [254:0]  io_input_payload_delay_2_stateElements_2;
  reg        [254:0]  io_input_payload_delay_2_stateElements_3;
  reg        [254:0]  io_input_payload_delay_2_stateElements_4;
  reg        [254:0]  io_input_payload_delay_2_stateElements_5;
  reg        [254:0]  io_input_payload_delay_2_stateElements_6;
  reg        [254:0]  io_input_payload_delay_2_stateElements_7;
  reg        [254:0]  io_input_payload_delay_2_stateElements_8;
  reg        [254:0]  io_input_payload_delay_2_stateElements_9;
  reg        [254:0]  io_input_payload_delay_2_stateElements_10;
  reg        [254:0]  io_input_payload_delay_2_stateElement;
  reg                 io_input_payload_delay_3_isFull;
  reg        [2:0]    io_input_payload_delay_3_fullRound;
  reg        [5:0]    io_input_payload_delay_3_partialRound;
  reg        [3:0]    io_input_payload_delay_3_stateIndex;
  reg        [3:0]    io_input_payload_delay_3_stateSize;
  reg        [7:0]    io_input_payload_delay_3_stateID;
  reg        [254:0]  io_input_payload_delay_3_stateElements_0;
  reg        [254:0]  io_input_payload_delay_3_stateElements_1;
  reg        [254:0]  io_input_payload_delay_3_stateElements_2;
  reg        [254:0]  io_input_payload_delay_3_stateElements_3;
  reg        [254:0]  io_input_payload_delay_3_stateElements_4;
  reg        [254:0]  io_input_payload_delay_3_stateElements_5;
  reg        [254:0]  io_input_payload_delay_3_stateElements_6;
  reg        [254:0]  io_input_payload_delay_3_stateElements_7;
  reg        [254:0]  io_input_payload_delay_3_stateElements_8;
  reg        [254:0]  io_input_payload_delay_3_stateElements_9;
  reg        [254:0]  io_input_payload_delay_3_stateElements_10;
  reg        [254:0]  io_input_payload_delay_3_stateElement;
  reg                 io_input_payload_delay_4_isFull;
  reg        [2:0]    io_input_payload_delay_4_fullRound;
  reg        [5:0]    io_input_payload_delay_4_partialRound;
  reg        [3:0]    io_input_payload_delay_4_stateIndex;
  reg        [3:0]    io_input_payload_delay_4_stateSize;
  reg        [7:0]    io_input_payload_delay_4_stateID;
  reg        [254:0]  io_input_payload_delay_4_stateElements_0;
  reg        [254:0]  io_input_payload_delay_4_stateElements_1;
  reg        [254:0]  io_input_payload_delay_4_stateElements_2;
  reg        [254:0]  io_input_payload_delay_4_stateElements_3;
  reg        [254:0]  io_input_payload_delay_4_stateElements_4;
  reg        [254:0]  io_input_payload_delay_4_stateElements_5;
  reg        [254:0]  io_input_payload_delay_4_stateElements_6;
  reg        [254:0]  io_input_payload_delay_4_stateElements_7;
  reg        [254:0]  io_input_payload_delay_4_stateElements_8;
  reg        [254:0]  io_input_payload_delay_4_stateElements_9;
  reg        [254:0]  io_input_payload_delay_4_stateElements_10;
  reg        [254:0]  io_input_payload_delay_4_stateElement;
  reg                 io_input_payload_delay_5_isFull;
  reg        [2:0]    io_input_payload_delay_5_fullRound;
  reg        [5:0]    io_input_payload_delay_5_partialRound;
  reg        [3:0]    io_input_payload_delay_5_stateIndex;
  reg        [3:0]    io_input_payload_delay_5_stateSize;
  reg        [7:0]    io_input_payload_delay_5_stateID;
  reg        [254:0]  io_input_payload_delay_5_stateElements_0;
  reg        [254:0]  io_input_payload_delay_5_stateElements_1;
  reg        [254:0]  io_input_payload_delay_5_stateElements_2;
  reg        [254:0]  io_input_payload_delay_5_stateElements_3;
  reg        [254:0]  io_input_payload_delay_5_stateElements_4;
  reg        [254:0]  io_input_payload_delay_5_stateElements_5;
  reg        [254:0]  io_input_payload_delay_5_stateElements_6;
  reg        [254:0]  io_input_payload_delay_5_stateElements_7;
  reg        [254:0]  io_input_payload_delay_5_stateElements_8;
  reg        [254:0]  io_input_payload_delay_5_stateElements_9;
  reg        [254:0]  io_input_payload_delay_5_stateElements_10;
  reg        [254:0]  io_input_payload_delay_5_stateElement;
  reg                 io_input_payload_delay_6_isFull;
  reg        [2:0]    io_input_payload_delay_6_fullRound;
  reg        [5:0]    io_input_payload_delay_6_partialRound;
  reg        [3:0]    io_input_payload_delay_6_stateIndex;
  reg        [3:0]    io_input_payload_delay_6_stateSize;
  reg        [7:0]    io_input_payload_delay_6_stateID;
  reg        [254:0]  io_input_payload_delay_6_stateElements_0;
  reg        [254:0]  io_input_payload_delay_6_stateElements_1;
  reg        [254:0]  io_input_payload_delay_6_stateElements_2;
  reg        [254:0]  io_input_payload_delay_6_stateElements_3;
  reg        [254:0]  io_input_payload_delay_6_stateElements_4;
  reg        [254:0]  io_input_payload_delay_6_stateElements_5;
  reg        [254:0]  io_input_payload_delay_6_stateElements_6;
  reg        [254:0]  io_input_payload_delay_6_stateElements_7;
  reg        [254:0]  io_input_payload_delay_6_stateElements_8;
  reg        [254:0]  io_input_payload_delay_6_stateElements_9;
  reg        [254:0]  io_input_payload_delay_6_stateElements_10;
  reg        [254:0]  io_input_payload_delay_6_stateElement;
  reg                 io_input_payload_delay_7_isFull;
  reg        [2:0]    io_input_payload_delay_7_fullRound;
  reg        [5:0]    io_input_payload_delay_7_partialRound;
  reg        [3:0]    io_input_payload_delay_7_stateIndex;
  reg        [3:0]    io_input_payload_delay_7_stateSize;
  reg        [7:0]    io_input_payload_delay_7_stateID;
  reg        [254:0]  io_input_payload_delay_7_stateElements_0;
  reg        [254:0]  io_input_payload_delay_7_stateElements_1;
  reg        [254:0]  io_input_payload_delay_7_stateElements_2;
  reg        [254:0]  io_input_payload_delay_7_stateElements_3;
  reg        [254:0]  io_input_payload_delay_7_stateElements_4;
  reg        [254:0]  io_input_payload_delay_7_stateElements_5;
  reg        [254:0]  io_input_payload_delay_7_stateElements_6;
  reg        [254:0]  io_input_payload_delay_7_stateElements_7;
  reg        [254:0]  io_input_payload_delay_7_stateElements_8;
  reg        [254:0]  io_input_payload_delay_7_stateElements_9;
  reg        [254:0]  io_input_payload_delay_7_stateElements_10;
  reg        [254:0]  io_input_payload_delay_7_stateElement;
  reg                 io_input_payload_delay_8_isFull;
  reg        [2:0]    io_input_payload_delay_8_fullRound;
  reg        [5:0]    io_input_payload_delay_8_partialRound;
  reg        [3:0]    io_input_payload_delay_8_stateIndex;
  reg        [3:0]    io_input_payload_delay_8_stateSize;
  reg        [7:0]    io_input_payload_delay_8_stateID;
  reg        [254:0]  io_input_payload_delay_8_stateElements_0;
  reg        [254:0]  io_input_payload_delay_8_stateElements_1;
  reg        [254:0]  io_input_payload_delay_8_stateElements_2;
  reg        [254:0]  io_input_payload_delay_8_stateElements_3;
  reg        [254:0]  io_input_payload_delay_8_stateElements_4;
  reg        [254:0]  io_input_payload_delay_8_stateElements_5;
  reg        [254:0]  io_input_payload_delay_8_stateElements_6;
  reg        [254:0]  io_input_payload_delay_8_stateElements_7;
  reg        [254:0]  io_input_payload_delay_8_stateElements_8;
  reg        [254:0]  io_input_payload_delay_8_stateElements_9;
  reg        [254:0]  io_input_payload_delay_8_stateElements_10;
  reg        [254:0]  io_input_payload_delay_8_stateElement;
  reg                 io_input_payload_delay_9_isFull;
  reg        [2:0]    io_input_payload_delay_9_fullRound;
  reg        [5:0]    io_input_payload_delay_9_partialRound;
  reg        [3:0]    io_input_payload_delay_9_stateIndex;
  reg        [3:0]    io_input_payload_delay_9_stateSize;
  reg        [7:0]    io_input_payload_delay_9_stateID;
  reg        [254:0]  io_input_payload_delay_9_stateElements_0;
  reg        [254:0]  io_input_payload_delay_9_stateElements_1;
  reg        [254:0]  io_input_payload_delay_9_stateElements_2;
  reg        [254:0]  io_input_payload_delay_9_stateElements_3;
  reg        [254:0]  io_input_payload_delay_9_stateElements_4;
  reg        [254:0]  io_input_payload_delay_9_stateElements_5;
  reg        [254:0]  io_input_payload_delay_9_stateElements_6;
  reg        [254:0]  io_input_payload_delay_9_stateElements_7;
  reg        [254:0]  io_input_payload_delay_9_stateElements_8;
  reg        [254:0]  io_input_payload_delay_9_stateElements_9;
  reg        [254:0]  io_input_payload_delay_9_stateElements_10;
  reg        [254:0]  io_input_payload_delay_9_stateElement;
  reg                 io_input_payload_delay_10_isFull;
  reg        [2:0]    io_input_payload_delay_10_fullRound;
  reg        [5:0]    io_input_payload_delay_10_partialRound;
  reg        [3:0]    io_input_payload_delay_10_stateIndex;
  reg        [3:0]    io_input_payload_delay_10_stateSize;
  reg        [7:0]    io_input_payload_delay_10_stateID;
  reg        [254:0]  io_input_payload_delay_10_stateElements_0;
  reg        [254:0]  io_input_payload_delay_10_stateElements_1;
  reg        [254:0]  io_input_payload_delay_10_stateElements_2;
  reg        [254:0]  io_input_payload_delay_10_stateElements_3;
  reg        [254:0]  io_input_payload_delay_10_stateElements_4;
  reg        [254:0]  io_input_payload_delay_10_stateElements_5;
  reg        [254:0]  io_input_payload_delay_10_stateElements_6;
  reg        [254:0]  io_input_payload_delay_10_stateElements_7;
  reg        [254:0]  io_input_payload_delay_10_stateElements_8;
  reg        [254:0]  io_input_payload_delay_10_stateElements_9;
  reg        [254:0]  io_input_payload_delay_10_stateElements_10;
  reg        [254:0]  io_input_payload_delay_10_stateElement;
  reg                 io_input_payload_delay_11_isFull;
  reg        [2:0]    io_input_payload_delay_11_fullRound;
  reg        [5:0]    io_input_payload_delay_11_partialRound;
  reg        [3:0]    io_input_payload_delay_11_stateIndex;
  reg        [3:0]    io_input_payload_delay_11_stateSize;
  reg        [7:0]    io_input_payload_delay_11_stateID;
  reg        [254:0]  io_input_payload_delay_11_stateElements_0;
  reg        [254:0]  io_input_payload_delay_11_stateElements_1;
  reg        [254:0]  io_input_payload_delay_11_stateElements_2;
  reg        [254:0]  io_input_payload_delay_11_stateElements_3;
  reg        [254:0]  io_input_payload_delay_11_stateElements_4;
  reg        [254:0]  io_input_payload_delay_11_stateElements_5;
  reg        [254:0]  io_input_payload_delay_11_stateElements_6;
  reg        [254:0]  io_input_payload_delay_11_stateElements_7;
  reg        [254:0]  io_input_payload_delay_11_stateElements_8;
  reg        [254:0]  io_input_payload_delay_11_stateElements_9;
  reg        [254:0]  io_input_payload_delay_11_stateElements_10;
  reg        [254:0]  io_input_payload_delay_11_stateElement;
  reg                 io_input_payload_delay_12_isFull;
  reg        [2:0]    io_input_payload_delay_12_fullRound;
  reg        [5:0]    io_input_payload_delay_12_partialRound;
  reg        [3:0]    io_input_payload_delay_12_stateIndex;
  reg        [3:0]    io_input_payload_delay_12_stateSize;
  reg        [7:0]    io_input_payload_delay_12_stateID;
  reg        [254:0]  io_input_payload_delay_12_stateElements_0;
  reg        [254:0]  io_input_payload_delay_12_stateElements_1;
  reg        [254:0]  io_input_payload_delay_12_stateElements_2;
  reg        [254:0]  io_input_payload_delay_12_stateElements_3;
  reg        [254:0]  io_input_payload_delay_12_stateElements_4;
  reg        [254:0]  io_input_payload_delay_12_stateElements_5;
  reg        [254:0]  io_input_payload_delay_12_stateElements_6;
  reg        [254:0]  io_input_payload_delay_12_stateElements_7;
  reg        [254:0]  io_input_payload_delay_12_stateElements_8;
  reg        [254:0]  io_input_payload_delay_12_stateElements_9;
  reg        [254:0]  io_input_payload_delay_12_stateElements_10;
  reg        [254:0]  io_input_payload_delay_12_stateElement;
  reg                 io_input_payload_delay_13_isFull;
  reg        [2:0]    io_input_payload_delay_13_fullRound;
  reg        [5:0]    io_input_payload_delay_13_partialRound;
  reg        [3:0]    io_input_payload_delay_13_stateIndex;
  reg        [3:0]    io_input_payload_delay_13_stateSize;
  reg        [7:0]    io_input_payload_delay_13_stateID;
  reg        [254:0]  io_input_payload_delay_13_stateElements_0;
  reg        [254:0]  io_input_payload_delay_13_stateElements_1;
  reg        [254:0]  io_input_payload_delay_13_stateElements_2;
  reg        [254:0]  io_input_payload_delay_13_stateElements_3;
  reg        [254:0]  io_input_payload_delay_13_stateElements_4;
  reg        [254:0]  io_input_payload_delay_13_stateElements_5;
  reg        [254:0]  io_input_payload_delay_13_stateElements_6;
  reg        [254:0]  io_input_payload_delay_13_stateElements_7;
  reg        [254:0]  io_input_payload_delay_13_stateElements_8;
  reg        [254:0]  io_input_payload_delay_13_stateElements_9;
  reg        [254:0]  io_input_payload_delay_13_stateElements_10;
  reg        [254:0]  io_input_payload_delay_13_stateElement;
  reg                 io_input_payload_delay_14_isFull;
  reg        [2:0]    io_input_payload_delay_14_fullRound;
  reg        [5:0]    io_input_payload_delay_14_partialRound;
  reg        [3:0]    io_input_payload_delay_14_stateIndex;
  reg        [3:0]    io_input_payload_delay_14_stateSize;
  reg        [7:0]    io_input_payload_delay_14_stateID;
  reg        [254:0]  io_input_payload_delay_14_stateElements_0;
  reg        [254:0]  io_input_payload_delay_14_stateElements_1;
  reg        [254:0]  io_input_payload_delay_14_stateElements_2;
  reg        [254:0]  io_input_payload_delay_14_stateElements_3;
  reg        [254:0]  io_input_payload_delay_14_stateElements_4;
  reg        [254:0]  io_input_payload_delay_14_stateElements_5;
  reg        [254:0]  io_input_payload_delay_14_stateElements_6;
  reg        [254:0]  io_input_payload_delay_14_stateElements_7;
  reg        [254:0]  io_input_payload_delay_14_stateElements_8;
  reg        [254:0]  io_input_payload_delay_14_stateElements_9;
  reg        [254:0]  io_input_payload_delay_14_stateElements_10;
  reg        [254:0]  io_input_payload_delay_14_stateElement;
  reg                 io_input_payload_delay_15_isFull;
  reg        [2:0]    io_input_payload_delay_15_fullRound;
  reg        [5:0]    io_input_payload_delay_15_partialRound;
  reg        [3:0]    io_input_payload_delay_15_stateIndex;
  reg        [3:0]    io_input_payload_delay_15_stateSize;
  reg        [7:0]    io_input_payload_delay_15_stateID;
  reg        [254:0]  io_input_payload_delay_15_stateElements_0;
  reg        [254:0]  io_input_payload_delay_15_stateElements_1;
  reg        [254:0]  io_input_payload_delay_15_stateElements_2;
  reg        [254:0]  io_input_payload_delay_15_stateElements_3;
  reg        [254:0]  io_input_payload_delay_15_stateElements_4;
  reg        [254:0]  io_input_payload_delay_15_stateElements_5;
  reg        [254:0]  io_input_payload_delay_15_stateElements_6;
  reg        [254:0]  io_input_payload_delay_15_stateElements_7;
  reg        [254:0]  io_input_payload_delay_15_stateElements_8;
  reg        [254:0]  io_input_payload_delay_15_stateElements_9;
  reg        [254:0]  io_input_payload_delay_15_stateElements_10;
  reg        [254:0]  io_input_payload_delay_15_stateElement;
  reg                 io_input_payload_delay_16_isFull;
  reg        [2:0]    io_input_payload_delay_16_fullRound;
  reg        [5:0]    io_input_payload_delay_16_partialRound;
  reg        [3:0]    io_input_payload_delay_16_stateIndex;
  reg        [3:0]    io_input_payload_delay_16_stateSize;
  reg        [7:0]    io_input_payload_delay_16_stateID;
  reg        [254:0]  io_input_payload_delay_16_stateElements_0;
  reg        [254:0]  io_input_payload_delay_16_stateElements_1;
  reg        [254:0]  io_input_payload_delay_16_stateElements_2;
  reg        [254:0]  io_input_payload_delay_16_stateElements_3;
  reg        [254:0]  io_input_payload_delay_16_stateElements_4;
  reg        [254:0]  io_input_payload_delay_16_stateElements_5;
  reg        [254:0]  io_input_payload_delay_16_stateElements_6;
  reg        [254:0]  io_input_payload_delay_16_stateElements_7;
  reg        [254:0]  io_input_payload_delay_16_stateElements_8;
  reg        [254:0]  io_input_payload_delay_16_stateElements_9;
  reg        [254:0]  io_input_payload_delay_16_stateElements_10;
  reg        [254:0]  io_input_payload_delay_16_stateElement;
  reg                 io_input_payload_delay_17_isFull;
  reg        [2:0]    io_input_payload_delay_17_fullRound;
  reg        [5:0]    io_input_payload_delay_17_partialRound;
  reg        [3:0]    io_input_payload_delay_17_stateIndex;
  reg        [3:0]    io_input_payload_delay_17_stateSize;
  reg        [7:0]    io_input_payload_delay_17_stateID;
  reg        [254:0]  io_input_payload_delay_17_stateElements_0;
  reg        [254:0]  io_input_payload_delay_17_stateElements_1;
  reg        [254:0]  io_input_payload_delay_17_stateElements_2;
  reg        [254:0]  io_input_payload_delay_17_stateElements_3;
  reg        [254:0]  io_input_payload_delay_17_stateElements_4;
  reg        [254:0]  io_input_payload_delay_17_stateElements_5;
  reg        [254:0]  io_input_payload_delay_17_stateElements_6;
  reg        [254:0]  io_input_payload_delay_17_stateElements_7;
  reg        [254:0]  io_input_payload_delay_17_stateElements_8;
  reg        [254:0]  io_input_payload_delay_17_stateElements_9;
  reg        [254:0]  io_input_payload_delay_17_stateElements_10;
  reg        [254:0]  io_input_payload_delay_17_stateElement;
  reg                 io_input_payload_delay_18_isFull;
  reg        [2:0]    io_input_payload_delay_18_fullRound;
  reg        [5:0]    io_input_payload_delay_18_partialRound;
  reg        [3:0]    io_input_payload_delay_18_stateIndex;
  reg        [3:0]    io_input_payload_delay_18_stateSize;
  reg        [7:0]    io_input_payload_delay_18_stateID;
  reg        [254:0]  io_input_payload_delay_18_stateElements_0;
  reg        [254:0]  io_input_payload_delay_18_stateElements_1;
  reg        [254:0]  io_input_payload_delay_18_stateElements_2;
  reg        [254:0]  io_input_payload_delay_18_stateElements_3;
  reg        [254:0]  io_input_payload_delay_18_stateElements_4;
  reg        [254:0]  io_input_payload_delay_18_stateElements_5;
  reg        [254:0]  io_input_payload_delay_18_stateElements_6;
  reg        [254:0]  io_input_payload_delay_18_stateElements_7;
  reg        [254:0]  io_input_payload_delay_18_stateElements_8;
  reg        [254:0]  io_input_payload_delay_18_stateElements_9;
  reg        [254:0]  io_input_payload_delay_18_stateElements_10;
  reg        [254:0]  io_input_payload_delay_18_stateElement;
  reg                 io_input_payload_delay_19_isFull;
  reg        [2:0]    io_input_payload_delay_19_fullRound;
  reg        [5:0]    io_input_payload_delay_19_partialRound;
  reg        [3:0]    io_input_payload_delay_19_stateIndex;
  reg        [3:0]    io_input_payload_delay_19_stateSize;
  reg        [7:0]    io_input_payload_delay_19_stateID;
  reg        [254:0]  io_input_payload_delay_19_stateElements_0;
  reg        [254:0]  io_input_payload_delay_19_stateElements_1;
  reg        [254:0]  io_input_payload_delay_19_stateElements_2;
  reg        [254:0]  io_input_payload_delay_19_stateElements_3;
  reg        [254:0]  io_input_payload_delay_19_stateElements_4;
  reg        [254:0]  io_input_payload_delay_19_stateElements_5;
  reg        [254:0]  io_input_payload_delay_19_stateElements_6;
  reg        [254:0]  io_input_payload_delay_19_stateElements_7;
  reg        [254:0]  io_input_payload_delay_19_stateElements_8;
  reg        [254:0]  io_input_payload_delay_19_stateElements_9;
  reg        [254:0]  io_input_payload_delay_19_stateElements_10;
  reg        [254:0]  io_input_payload_delay_19_stateElement;
  reg                 io_input_payload_delay_20_isFull;
  reg        [2:0]    io_input_payload_delay_20_fullRound;
  reg        [5:0]    io_input_payload_delay_20_partialRound;
  reg        [3:0]    io_input_payload_delay_20_stateIndex;
  reg        [3:0]    io_input_payload_delay_20_stateSize;
  reg        [7:0]    io_input_payload_delay_20_stateID;
  reg        [254:0]  io_input_payload_delay_20_stateElements_0;
  reg        [254:0]  io_input_payload_delay_20_stateElements_1;
  reg        [254:0]  io_input_payload_delay_20_stateElements_2;
  reg        [254:0]  io_input_payload_delay_20_stateElements_3;
  reg        [254:0]  io_input_payload_delay_20_stateElements_4;
  reg        [254:0]  io_input_payload_delay_20_stateElements_5;
  reg        [254:0]  io_input_payload_delay_20_stateElements_6;
  reg        [254:0]  io_input_payload_delay_20_stateElements_7;
  reg        [254:0]  io_input_payload_delay_20_stateElements_8;
  reg        [254:0]  io_input_payload_delay_20_stateElements_9;
  reg        [254:0]  io_input_payload_delay_20_stateElements_10;
  reg        [254:0]  io_input_payload_delay_20_stateElement;
  reg                 io_input_payload_delay_21_isFull;
  reg        [2:0]    io_input_payload_delay_21_fullRound;
  reg        [5:0]    io_input_payload_delay_21_partialRound;
  reg        [3:0]    io_input_payload_delay_21_stateIndex;
  reg        [3:0]    io_input_payload_delay_21_stateSize;
  reg        [7:0]    io_input_payload_delay_21_stateID;
  reg        [254:0]  io_input_payload_delay_21_stateElements_0;
  reg        [254:0]  io_input_payload_delay_21_stateElements_1;
  reg        [254:0]  io_input_payload_delay_21_stateElements_2;
  reg        [254:0]  io_input_payload_delay_21_stateElements_3;
  reg        [254:0]  io_input_payload_delay_21_stateElements_4;
  reg        [254:0]  io_input_payload_delay_21_stateElements_5;
  reg        [254:0]  io_input_payload_delay_21_stateElements_6;
  reg        [254:0]  io_input_payload_delay_21_stateElements_7;
  reg        [254:0]  io_input_payload_delay_21_stateElements_8;
  reg        [254:0]  io_input_payload_delay_21_stateElements_9;
  reg        [254:0]  io_input_payload_delay_21_stateElements_10;
  reg        [254:0]  io_input_payload_delay_21_stateElement;
  reg                 io_input_payload_delay_22_isFull;
  reg        [2:0]    io_input_payload_delay_22_fullRound;
  reg        [5:0]    io_input_payload_delay_22_partialRound;
  reg        [3:0]    io_input_payload_delay_22_stateIndex;
  reg        [3:0]    io_input_payload_delay_22_stateSize;
  reg        [7:0]    io_input_payload_delay_22_stateID;
  reg        [254:0]  io_input_payload_delay_22_stateElements_0;
  reg        [254:0]  io_input_payload_delay_22_stateElements_1;
  reg        [254:0]  io_input_payload_delay_22_stateElements_2;
  reg        [254:0]  io_input_payload_delay_22_stateElements_3;
  reg        [254:0]  io_input_payload_delay_22_stateElements_4;
  reg        [254:0]  io_input_payload_delay_22_stateElements_5;
  reg        [254:0]  io_input_payload_delay_22_stateElements_6;
  reg        [254:0]  io_input_payload_delay_22_stateElements_7;
  reg        [254:0]  io_input_payload_delay_22_stateElements_8;
  reg        [254:0]  io_input_payload_delay_22_stateElements_9;
  reg        [254:0]  io_input_payload_delay_22_stateElements_10;
  reg        [254:0]  io_input_payload_delay_22_stateElement;
  reg                 io_input_payload_delay_23_isFull;
  reg        [2:0]    io_input_payload_delay_23_fullRound;
  reg        [5:0]    io_input_payload_delay_23_partialRound;
  reg        [3:0]    io_input_payload_delay_23_stateIndex;
  reg        [3:0]    io_input_payload_delay_23_stateSize;
  reg        [7:0]    io_input_payload_delay_23_stateID;
  reg        [254:0]  io_input_payload_delay_23_stateElements_0;
  reg        [254:0]  io_input_payload_delay_23_stateElements_1;
  reg        [254:0]  io_input_payload_delay_23_stateElements_2;
  reg        [254:0]  io_input_payload_delay_23_stateElements_3;
  reg        [254:0]  io_input_payload_delay_23_stateElements_4;
  reg        [254:0]  io_input_payload_delay_23_stateElements_5;
  reg        [254:0]  io_input_payload_delay_23_stateElements_6;
  reg        [254:0]  io_input_payload_delay_23_stateElements_7;
  reg        [254:0]  io_input_payload_delay_23_stateElements_8;
  reg        [254:0]  io_input_payload_delay_23_stateElements_9;
  reg        [254:0]  io_input_payload_delay_23_stateElements_10;
  reg        [254:0]  io_input_payload_delay_23_stateElement;
  reg                 io_input_payload_delay_24_isFull;
  reg        [2:0]    io_input_payload_delay_24_fullRound;
  reg        [5:0]    io_input_payload_delay_24_partialRound;
  reg        [3:0]    io_input_payload_delay_24_stateIndex;
  reg        [3:0]    io_input_payload_delay_24_stateSize;
  reg        [7:0]    io_input_payload_delay_24_stateID;
  reg        [254:0]  io_input_payload_delay_24_stateElements_0;
  reg        [254:0]  io_input_payload_delay_24_stateElements_1;
  reg        [254:0]  io_input_payload_delay_24_stateElements_2;
  reg        [254:0]  io_input_payload_delay_24_stateElements_3;
  reg        [254:0]  io_input_payload_delay_24_stateElements_4;
  reg        [254:0]  io_input_payload_delay_24_stateElements_5;
  reg        [254:0]  io_input_payload_delay_24_stateElements_6;
  reg        [254:0]  io_input_payload_delay_24_stateElements_7;
  reg        [254:0]  io_input_payload_delay_24_stateElements_8;
  reg        [254:0]  io_input_payload_delay_24_stateElements_9;
  reg        [254:0]  io_input_payload_delay_24_stateElements_10;
  reg        [254:0]  io_input_payload_delay_24_stateElement;
  reg                 io_input_payload_delay_25_isFull;
  reg        [2:0]    io_input_payload_delay_25_fullRound;
  reg        [5:0]    io_input_payload_delay_25_partialRound;
  reg        [3:0]    io_input_payload_delay_25_stateIndex;
  reg        [3:0]    io_input_payload_delay_25_stateSize;
  reg        [7:0]    io_input_payload_delay_25_stateID;
  reg        [254:0]  io_input_payload_delay_25_stateElements_0;
  reg        [254:0]  io_input_payload_delay_25_stateElements_1;
  reg        [254:0]  io_input_payload_delay_25_stateElements_2;
  reg        [254:0]  io_input_payload_delay_25_stateElements_3;
  reg        [254:0]  io_input_payload_delay_25_stateElements_4;
  reg        [254:0]  io_input_payload_delay_25_stateElements_5;
  reg        [254:0]  io_input_payload_delay_25_stateElements_6;
  reg        [254:0]  io_input_payload_delay_25_stateElements_7;
  reg        [254:0]  io_input_payload_delay_25_stateElements_8;
  reg        [254:0]  io_input_payload_delay_25_stateElements_9;
  reg        [254:0]  io_input_payload_delay_25_stateElements_10;
  reg        [254:0]  io_input_payload_delay_25_stateElement;
  reg                 io_input_payload_delay_26_isFull;
  reg        [2:0]    io_input_payload_delay_26_fullRound;
  reg        [5:0]    io_input_payload_delay_26_partialRound;
  reg        [3:0]    io_input_payload_delay_26_stateIndex;
  reg        [3:0]    io_input_payload_delay_26_stateSize;
  reg        [7:0]    io_input_payload_delay_26_stateID;
  reg        [254:0]  io_input_payload_delay_26_stateElements_0;
  reg        [254:0]  io_input_payload_delay_26_stateElements_1;
  reg        [254:0]  io_input_payload_delay_26_stateElements_2;
  reg        [254:0]  io_input_payload_delay_26_stateElements_3;
  reg        [254:0]  io_input_payload_delay_26_stateElements_4;
  reg        [254:0]  io_input_payload_delay_26_stateElements_5;
  reg        [254:0]  io_input_payload_delay_26_stateElements_6;
  reg        [254:0]  io_input_payload_delay_26_stateElements_7;
  reg        [254:0]  io_input_payload_delay_26_stateElements_8;
  reg        [254:0]  io_input_payload_delay_26_stateElements_9;
  reg        [254:0]  io_input_payload_delay_26_stateElements_10;
  reg        [254:0]  io_input_payload_delay_26_stateElement;
  reg                 io_input_payload_delay_27_isFull;
  reg        [2:0]    io_input_payload_delay_27_fullRound;
  reg        [5:0]    io_input_payload_delay_27_partialRound;
  reg        [3:0]    io_input_payload_delay_27_stateIndex;
  reg        [3:0]    io_input_payload_delay_27_stateSize;
  reg        [7:0]    io_input_payload_delay_27_stateID;
  reg        [254:0]  io_input_payload_delay_27_stateElements_0;
  reg        [254:0]  io_input_payload_delay_27_stateElements_1;
  reg        [254:0]  io_input_payload_delay_27_stateElements_2;
  reg        [254:0]  io_input_payload_delay_27_stateElements_3;
  reg        [254:0]  io_input_payload_delay_27_stateElements_4;
  reg        [254:0]  io_input_payload_delay_27_stateElements_5;
  reg        [254:0]  io_input_payload_delay_27_stateElements_6;
  reg        [254:0]  io_input_payload_delay_27_stateElements_7;
  reg        [254:0]  io_input_payload_delay_27_stateElements_8;
  reg        [254:0]  io_input_payload_delay_27_stateElements_9;
  reg        [254:0]  io_input_payload_delay_27_stateElements_10;
  reg        [254:0]  io_input_payload_delay_27_stateElement;
  reg                 io_input_payload_delay_28_isFull;
  reg        [2:0]    io_input_payload_delay_28_fullRound;
  reg        [5:0]    io_input_payload_delay_28_partialRound;
  reg        [3:0]    io_input_payload_delay_28_stateIndex;
  reg        [3:0]    io_input_payload_delay_28_stateSize;
  reg        [7:0]    io_input_payload_delay_28_stateID;
  reg        [254:0]  io_input_payload_delay_28_stateElements_0;
  reg        [254:0]  io_input_payload_delay_28_stateElements_1;
  reg        [254:0]  io_input_payload_delay_28_stateElements_2;
  reg        [254:0]  io_input_payload_delay_28_stateElements_3;
  reg        [254:0]  io_input_payload_delay_28_stateElements_4;
  reg        [254:0]  io_input_payload_delay_28_stateElements_5;
  reg        [254:0]  io_input_payload_delay_28_stateElements_6;
  reg        [254:0]  io_input_payload_delay_28_stateElements_7;
  reg        [254:0]  io_input_payload_delay_28_stateElements_8;
  reg        [254:0]  io_input_payload_delay_28_stateElements_9;
  reg        [254:0]  io_input_payload_delay_28_stateElements_10;
  reg        [254:0]  io_input_payload_delay_28_stateElement;
  reg                 io_input_payload_delay_29_isFull;
  reg        [2:0]    io_input_payload_delay_29_fullRound;
  reg        [5:0]    io_input_payload_delay_29_partialRound;
  reg        [3:0]    io_input_payload_delay_29_stateIndex;
  reg        [3:0]    io_input_payload_delay_29_stateSize;
  reg        [7:0]    io_input_payload_delay_29_stateID;
  reg        [254:0]  io_input_payload_delay_29_stateElements_0;
  reg        [254:0]  io_input_payload_delay_29_stateElements_1;
  reg        [254:0]  io_input_payload_delay_29_stateElements_2;
  reg        [254:0]  io_input_payload_delay_29_stateElements_3;
  reg        [254:0]  io_input_payload_delay_29_stateElements_4;
  reg        [254:0]  io_input_payload_delay_29_stateElements_5;
  reg        [254:0]  io_input_payload_delay_29_stateElements_6;
  reg        [254:0]  io_input_payload_delay_29_stateElements_7;
  reg        [254:0]  io_input_payload_delay_29_stateElements_8;
  reg        [254:0]  io_input_payload_delay_29_stateElements_9;
  reg        [254:0]  io_input_payload_delay_29_stateElements_10;
  reg        [254:0]  io_input_payload_delay_29_stateElement;
  reg                 io_input_payload_delay_30_isFull;
  reg        [2:0]    io_input_payload_delay_30_fullRound;
  reg        [5:0]    io_input_payload_delay_30_partialRound;
  reg        [3:0]    io_input_payload_delay_30_stateIndex;
  reg        [3:0]    io_input_payload_delay_30_stateSize;
  reg        [7:0]    io_input_payload_delay_30_stateID;
  reg        [254:0]  io_input_payload_delay_30_stateElements_0;
  reg        [254:0]  io_input_payload_delay_30_stateElements_1;
  reg        [254:0]  io_input_payload_delay_30_stateElements_2;
  reg        [254:0]  io_input_payload_delay_30_stateElements_3;
  reg        [254:0]  io_input_payload_delay_30_stateElements_4;
  reg        [254:0]  io_input_payload_delay_30_stateElements_5;
  reg        [254:0]  io_input_payload_delay_30_stateElements_6;
  reg        [254:0]  io_input_payload_delay_30_stateElements_7;
  reg        [254:0]  io_input_payload_delay_30_stateElements_8;
  reg        [254:0]  io_input_payload_delay_30_stateElements_9;
  reg        [254:0]  io_input_payload_delay_30_stateElements_10;
  reg        [254:0]  io_input_payload_delay_30_stateElement;
  reg                 io_input_payload_delay_31_isFull;
  reg        [2:0]    io_input_payload_delay_31_fullRound;
  reg        [5:0]    io_input_payload_delay_31_partialRound;
  reg        [3:0]    io_input_payload_delay_31_stateIndex;
  reg        [3:0]    io_input_payload_delay_31_stateSize;
  reg        [7:0]    io_input_payload_delay_31_stateID;
  reg        [254:0]  io_input_payload_delay_31_stateElements_0;
  reg        [254:0]  io_input_payload_delay_31_stateElements_1;
  reg        [254:0]  io_input_payload_delay_31_stateElements_2;
  reg        [254:0]  io_input_payload_delay_31_stateElements_3;
  reg        [254:0]  io_input_payload_delay_31_stateElements_4;
  reg        [254:0]  io_input_payload_delay_31_stateElements_5;
  reg        [254:0]  io_input_payload_delay_31_stateElements_6;
  reg        [254:0]  io_input_payload_delay_31_stateElements_7;
  reg        [254:0]  io_input_payload_delay_31_stateElements_8;
  reg        [254:0]  io_input_payload_delay_31_stateElements_9;
  reg        [254:0]  io_input_payload_delay_31_stateElements_10;
  reg        [254:0]  io_input_payload_delay_31_stateElement;
  reg                 io_input_payload_delay_32_isFull;
  reg        [2:0]    io_input_payload_delay_32_fullRound;
  reg        [5:0]    io_input_payload_delay_32_partialRound;
  reg        [3:0]    io_input_payload_delay_32_stateIndex;
  reg        [3:0]    io_input_payload_delay_32_stateSize;
  reg        [7:0]    io_input_payload_delay_32_stateID;
  reg        [254:0]  io_input_payload_delay_32_stateElements_0;
  reg        [254:0]  io_input_payload_delay_32_stateElements_1;
  reg        [254:0]  io_input_payload_delay_32_stateElements_2;
  reg        [254:0]  io_input_payload_delay_32_stateElements_3;
  reg        [254:0]  io_input_payload_delay_32_stateElements_4;
  reg        [254:0]  io_input_payload_delay_32_stateElements_5;
  reg        [254:0]  io_input_payload_delay_32_stateElements_6;
  reg        [254:0]  io_input_payload_delay_32_stateElements_7;
  reg        [254:0]  io_input_payload_delay_32_stateElements_8;
  reg        [254:0]  io_input_payload_delay_32_stateElements_9;
  reg        [254:0]  io_input_payload_delay_32_stateElements_10;
  reg        [254:0]  io_input_payload_delay_32_stateElement;
  reg                 io_input_payload_delay_33_isFull;
  reg        [2:0]    io_input_payload_delay_33_fullRound;
  reg        [5:0]    io_input_payload_delay_33_partialRound;
  reg        [3:0]    io_input_payload_delay_33_stateIndex;
  reg        [3:0]    io_input_payload_delay_33_stateSize;
  reg        [7:0]    io_input_payload_delay_33_stateID;
  reg        [254:0]  io_input_payload_delay_33_stateElements_0;
  reg        [254:0]  io_input_payload_delay_33_stateElements_1;
  reg        [254:0]  io_input_payload_delay_33_stateElements_2;
  reg        [254:0]  io_input_payload_delay_33_stateElements_3;
  reg        [254:0]  io_input_payload_delay_33_stateElements_4;
  reg        [254:0]  io_input_payload_delay_33_stateElements_5;
  reg        [254:0]  io_input_payload_delay_33_stateElements_6;
  reg        [254:0]  io_input_payload_delay_33_stateElements_7;
  reg        [254:0]  io_input_payload_delay_33_stateElements_8;
  reg        [254:0]  io_input_payload_delay_33_stateElements_9;
  reg        [254:0]  io_input_payload_delay_33_stateElements_10;
  reg        [254:0]  io_input_payload_delay_33_stateElement;
  reg                 io_input_payload_delay_34_isFull;
  reg        [2:0]    io_input_payload_delay_34_fullRound;
  reg        [5:0]    io_input_payload_delay_34_partialRound;
  reg        [3:0]    io_input_payload_delay_34_stateIndex;
  reg        [3:0]    io_input_payload_delay_34_stateSize;
  reg        [7:0]    io_input_payload_delay_34_stateID;
  reg        [254:0]  io_input_payload_delay_34_stateElements_0;
  reg        [254:0]  io_input_payload_delay_34_stateElements_1;
  reg        [254:0]  io_input_payload_delay_34_stateElements_2;
  reg        [254:0]  io_input_payload_delay_34_stateElements_3;
  reg        [254:0]  io_input_payload_delay_34_stateElements_4;
  reg        [254:0]  io_input_payload_delay_34_stateElements_5;
  reg        [254:0]  io_input_payload_delay_34_stateElements_6;
  reg        [254:0]  io_input_payload_delay_34_stateElements_7;
  reg        [254:0]  io_input_payload_delay_34_stateElements_8;
  reg        [254:0]  io_input_payload_delay_34_stateElements_9;
  reg        [254:0]  io_input_payload_delay_34_stateElements_10;
  reg        [254:0]  io_input_payload_delay_34_stateElement;
  reg                 io_input_payload_delay_35_isFull;
  reg        [2:0]    io_input_payload_delay_35_fullRound;
  reg        [5:0]    io_input_payload_delay_35_partialRound;
  reg        [3:0]    io_input_payload_delay_35_stateIndex;
  reg        [3:0]    io_input_payload_delay_35_stateSize;
  reg        [7:0]    io_input_payload_delay_35_stateID;
  reg        [254:0]  io_input_payload_delay_35_stateElements_0;
  reg        [254:0]  io_input_payload_delay_35_stateElements_1;
  reg        [254:0]  io_input_payload_delay_35_stateElements_2;
  reg        [254:0]  io_input_payload_delay_35_stateElements_3;
  reg        [254:0]  io_input_payload_delay_35_stateElements_4;
  reg        [254:0]  io_input_payload_delay_35_stateElements_5;
  reg        [254:0]  io_input_payload_delay_35_stateElements_6;
  reg        [254:0]  io_input_payload_delay_35_stateElements_7;
  reg        [254:0]  io_input_payload_delay_35_stateElements_8;
  reg        [254:0]  io_input_payload_delay_35_stateElements_9;
  reg        [254:0]  io_input_payload_delay_35_stateElements_10;
  reg        [254:0]  io_input_payload_delay_35_stateElement;
  reg                 io_input_payload_delay_36_isFull;
  reg        [2:0]    io_input_payload_delay_36_fullRound;
  reg        [5:0]    io_input_payload_delay_36_partialRound;
  reg        [3:0]    io_input_payload_delay_36_stateIndex;
  reg        [3:0]    io_input_payload_delay_36_stateSize;
  reg        [7:0]    io_input_payload_delay_36_stateID;
  reg        [254:0]  io_input_payload_delay_36_stateElements_0;
  reg        [254:0]  io_input_payload_delay_36_stateElements_1;
  reg        [254:0]  io_input_payload_delay_36_stateElements_2;
  reg        [254:0]  io_input_payload_delay_36_stateElements_3;
  reg        [254:0]  io_input_payload_delay_36_stateElements_4;
  reg        [254:0]  io_input_payload_delay_36_stateElements_5;
  reg        [254:0]  io_input_payload_delay_36_stateElements_6;
  reg        [254:0]  io_input_payload_delay_36_stateElements_7;
  reg        [254:0]  io_input_payload_delay_36_stateElements_8;
  reg        [254:0]  io_input_payload_delay_36_stateElements_9;
  reg        [254:0]  io_input_payload_delay_36_stateElements_10;
  reg        [254:0]  io_input_payload_delay_36_stateElement;
  reg                 io_input_payload_delay_37_isFull;
  reg        [2:0]    io_input_payload_delay_37_fullRound;
  reg        [5:0]    io_input_payload_delay_37_partialRound;
  reg        [3:0]    io_input_payload_delay_37_stateIndex;
  reg        [3:0]    io_input_payload_delay_37_stateSize;
  reg        [7:0]    io_input_payload_delay_37_stateID;
  reg        [254:0]  io_input_payload_delay_37_stateElements_0;
  reg        [254:0]  io_input_payload_delay_37_stateElements_1;
  reg        [254:0]  io_input_payload_delay_37_stateElements_2;
  reg        [254:0]  io_input_payload_delay_37_stateElements_3;
  reg        [254:0]  io_input_payload_delay_37_stateElements_4;
  reg        [254:0]  io_input_payload_delay_37_stateElements_5;
  reg        [254:0]  io_input_payload_delay_37_stateElements_6;
  reg        [254:0]  io_input_payload_delay_37_stateElements_7;
  reg        [254:0]  io_input_payload_delay_37_stateElements_8;
  reg        [254:0]  io_input_payload_delay_37_stateElements_9;
  reg        [254:0]  io_input_payload_delay_37_stateElements_10;
  reg        [254:0]  io_input_payload_delay_37_stateElement;
  reg                 io_input_payload_delay_38_isFull;
  reg        [2:0]    io_input_payload_delay_38_fullRound;
  reg        [5:0]    io_input_payload_delay_38_partialRound;
  reg        [3:0]    io_input_payload_delay_38_stateIndex;
  reg        [3:0]    io_input_payload_delay_38_stateSize;
  reg        [7:0]    io_input_payload_delay_38_stateID;
  reg        [254:0]  io_input_payload_delay_38_stateElements_0;
  reg        [254:0]  io_input_payload_delay_38_stateElements_1;
  reg        [254:0]  io_input_payload_delay_38_stateElements_2;
  reg        [254:0]  io_input_payload_delay_38_stateElements_3;
  reg        [254:0]  io_input_payload_delay_38_stateElements_4;
  reg        [254:0]  io_input_payload_delay_38_stateElements_5;
  reg        [254:0]  io_input_payload_delay_38_stateElements_6;
  reg        [254:0]  io_input_payload_delay_38_stateElements_7;
  reg        [254:0]  io_input_payload_delay_38_stateElements_8;
  reg        [254:0]  io_input_payload_delay_38_stateElements_9;
  reg        [254:0]  io_input_payload_delay_38_stateElements_10;
  reg        [254:0]  io_input_payload_delay_38_stateElement;
  reg                 io_input_payload_delay_39_isFull;
  reg        [2:0]    io_input_payload_delay_39_fullRound;
  reg        [5:0]    io_input_payload_delay_39_partialRound;
  reg        [3:0]    io_input_payload_delay_39_stateIndex;
  reg        [3:0]    io_input_payload_delay_39_stateSize;
  reg        [7:0]    io_input_payload_delay_39_stateID;
  reg        [254:0]  io_input_payload_delay_39_stateElements_0;
  reg        [254:0]  io_input_payload_delay_39_stateElements_1;
  reg        [254:0]  io_input_payload_delay_39_stateElements_2;
  reg        [254:0]  io_input_payload_delay_39_stateElements_3;
  reg        [254:0]  io_input_payload_delay_39_stateElements_4;
  reg        [254:0]  io_input_payload_delay_39_stateElements_5;
  reg        [254:0]  io_input_payload_delay_39_stateElements_6;
  reg        [254:0]  io_input_payload_delay_39_stateElements_7;
  reg        [254:0]  io_input_payload_delay_39_stateElements_8;
  reg        [254:0]  io_input_payload_delay_39_stateElements_9;
  reg        [254:0]  io_input_payload_delay_39_stateElements_10;
  reg        [254:0]  io_input_payload_delay_39_stateElement;
  reg                 io_input_payload_delay_40_isFull;
  reg        [2:0]    io_input_payload_delay_40_fullRound;
  reg        [5:0]    io_input_payload_delay_40_partialRound;
  reg        [3:0]    io_input_payload_delay_40_stateIndex;
  reg        [3:0]    io_input_payload_delay_40_stateSize;
  reg        [7:0]    io_input_payload_delay_40_stateID;
  reg        [254:0]  io_input_payload_delay_40_stateElements_0;
  reg        [254:0]  io_input_payload_delay_40_stateElements_1;
  reg        [254:0]  io_input_payload_delay_40_stateElements_2;
  reg        [254:0]  io_input_payload_delay_40_stateElements_3;
  reg        [254:0]  io_input_payload_delay_40_stateElements_4;
  reg        [254:0]  io_input_payload_delay_40_stateElements_5;
  reg        [254:0]  io_input_payload_delay_40_stateElements_6;
  reg        [254:0]  io_input_payload_delay_40_stateElements_7;
  reg        [254:0]  io_input_payload_delay_40_stateElements_8;
  reg        [254:0]  io_input_payload_delay_40_stateElements_9;
  reg        [254:0]  io_input_payload_delay_40_stateElements_10;
  reg        [254:0]  io_input_payload_delay_40_stateElement;
  reg                 io_input_payload_delay_41_isFull;
  reg        [2:0]    io_input_payload_delay_41_fullRound;
  reg        [5:0]    io_input_payload_delay_41_partialRound;
  reg        [3:0]    io_input_payload_delay_41_stateIndex;
  reg        [3:0]    io_input_payload_delay_41_stateSize;
  reg        [7:0]    io_input_payload_delay_41_stateID;
  reg        [254:0]  io_input_payload_delay_41_stateElements_0;
  reg        [254:0]  io_input_payload_delay_41_stateElements_1;
  reg        [254:0]  io_input_payload_delay_41_stateElements_2;
  reg        [254:0]  io_input_payload_delay_41_stateElements_3;
  reg        [254:0]  io_input_payload_delay_41_stateElements_4;
  reg        [254:0]  io_input_payload_delay_41_stateElements_5;
  reg        [254:0]  io_input_payload_delay_41_stateElements_6;
  reg        [254:0]  io_input_payload_delay_41_stateElements_7;
  reg        [254:0]  io_input_payload_delay_41_stateElements_8;
  reg        [254:0]  io_input_payload_delay_41_stateElements_9;
  reg        [254:0]  io_input_payload_delay_41_stateElements_10;
  reg        [254:0]  io_input_payload_delay_41_stateElement;
  reg                 io_input_payload_delay_42_isFull;
  reg        [2:0]    io_input_payload_delay_42_fullRound;
  reg        [5:0]    io_input_payload_delay_42_partialRound;
  reg        [3:0]    io_input_payload_delay_42_stateIndex;
  reg        [3:0]    io_input_payload_delay_42_stateSize;
  reg        [7:0]    io_input_payload_delay_42_stateID;
  reg        [254:0]  io_input_payload_delay_42_stateElements_0;
  reg        [254:0]  io_input_payload_delay_42_stateElements_1;
  reg        [254:0]  io_input_payload_delay_42_stateElements_2;
  reg        [254:0]  io_input_payload_delay_42_stateElements_3;
  reg        [254:0]  io_input_payload_delay_42_stateElements_4;
  reg        [254:0]  io_input_payload_delay_42_stateElements_5;
  reg        [254:0]  io_input_payload_delay_42_stateElements_6;
  reg        [254:0]  io_input_payload_delay_42_stateElements_7;
  reg        [254:0]  io_input_payload_delay_42_stateElements_8;
  reg        [254:0]  io_input_payload_delay_42_stateElements_9;
  reg        [254:0]  io_input_payload_delay_42_stateElements_10;
  reg        [254:0]  io_input_payload_delay_42_stateElement;
  reg                 io_input_payload_delay_43_isFull;
  reg        [2:0]    io_input_payload_delay_43_fullRound;
  reg        [5:0]    io_input_payload_delay_43_partialRound;
  reg        [3:0]    io_input_payload_delay_43_stateIndex;
  reg        [3:0]    io_input_payload_delay_43_stateSize;
  reg        [7:0]    io_input_payload_delay_43_stateID;
  reg        [254:0]  io_input_payload_delay_43_stateElements_0;
  reg        [254:0]  io_input_payload_delay_43_stateElements_1;
  reg        [254:0]  io_input_payload_delay_43_stateElements_2;
  reg        [254:0]  io_input_payload_delay_43_stateElements_3;
  reg        [254:0]  io_input_payload_delay_43_stateElements_4;
  reg        [254:0]  io_input_payload_delay_43_stateElements_5;
  reg        [254:0]  io_input_payload_delay_43_stateElements_6;
  reg        [254:0]  io_input_payload_delay_43_stateElements_7;
  reg        [254:0]  io_input_payload_delay_43_stateElements_8;
  reg        [254:0]  io_input_payload_delay_43_stateElements_9;
  reg        [254:0]  io_input_payload_delay_43_stateElements_10;
  reg        [254:0]  io_input_payload_delay_43_stateElement;
  reg                 io_input_payload_delay_44_isFull;
  reg        [2:0]    io_input_payload_delay_44_fullRound;
  reg        [5:0]    io_input_payload_delay_44_partialRound;
  reg        [3:0]    io_input_payload_delay_44_stateIndex;
  reg        [3:0]    io_input_payload_delay_44_stateSize;
  reg        [7:0]    io_input_payload_delay_44_stateID;
  reg        [254:0]  io_input_payload_delay_44_stateElements_0;
  reg        [254:0]  io_input_payload_delay_44_stateElements_1;
  reg        [254:0]  io_input_payload_delay_44_stateElements_2;
  reg        [254:0]  io_input_payload_delay_44_stateElements_3;
  reg        [254:0]  io_input_payload_delay_44_stateElements_4;
  reg        [254:0]  io_input_payload_delay_44_stateElements_5;
  reg        [254:0]  io_input_payload_delay_44_stateElements_6;
  reg        [254:0]  io_input_payload_delay_44_stateElements_7;
  reg        [254:0]  io_input_payload_delay_44_stateElements_8;
  reg        [254:0]  io_input_payload_delay_44_stateElements_9;
  reg        [254:0]  io_input_payload_delay_44_stateElements_10;
  reg        [254:0]  io_input_payload_delay_44_stateElement;
  reg                 io_input_payload_delay_45_isFull;
  reg        [2:0]    io_input_payload_delay_45_fullRound;
  reg        [5:0]    io_input_payload_delay_45_partialRound;
  reg        [3:0]    io_input_payload_delay_45_stateIndex;
  reg        [3:0]    io_input_payload_delay_45_stateSize;
  reg        [7:0]    io_input_payload_delay_45_stateID;
  reg        [254:0]  io_input_payload_delay_45_stateElements_0;
  reg        [254:0]  io_input_payload_delay_45_stateElements_1;
  reg        [254:0]  io_input_payload_delay_45_stateElements_2;
  reg        [254:0]  io_input_payload_delay_45_stateElements_3;
  reg        [254:0]  io_input_payload_delay_45_stateElements_4;
  reg        [254:0]  io_input_payload_delay_45_stateElements_5;
  reg        [254:0]  io_input_payload_delay_45_stateElements_6;
  reg        [254:0]  io_input_payload_delay_45_stateElements_7;
  reg        [254:0]  io_input_payload_delay_45_stateElements_8;
  reg        [254:0]  io_input_payload_delay_45_stateElements_9;
  reg        [254:0]  io_input_payload_delay_45_stateElements_10;
  reg        [254:0]  io_input_payload_delay_45_stateElement;
  reg                 io_input_payload_delay_46_isFull;
  reg        [2:0]    io_input_payload_delay_46_fullRound;
  reg        [5:0]    io_input_payload_delay_46_partialRound;
  reg        [3:0]    io_input_payload_delay_46_stateIndex;
  reg        [3:0]    io_input_payload_delay_46_stateSize;
  reg        [7:0]    io_input_payload_delay_46_stateID;
  reg        [254:0]  io_input_payload_delay_46_stateElements_0;
  reg        [254:0]  io_input_payload_delay_46_stateElements_1;
  reg        [254:0]  io_input_payload_delay_46_stateElements_2;
  reg        [254:0]  io_input_payload_delay_46_stateElements_3;
  reg        [254:0]  io_input_payload_delay_46_stateElements_4;
  reg        [254:0]  io_input_payload_delay_46_stateElements_5;
  reg        [254:0]  io_input_payload_delay_46_stateElements_6;
  reg        [254:0]  io_input_payload_delay_46_stateElements_7;
  reg        [254:0]  io_input_payload_delay_46_stateElements_8;
  reg        [254:0]  io_input_payload_delay_46_stateElements_9;
  reg        [254:0]  io_input_payload_delay_46_stateElements_10;
  reg        [254:0]  io_input_payload_delay_46_stateElement;
  reg                 io_input_payload_delay_47_isFull;
  reg        [2:0]    io_input_payload_delay_47_fullRound;
  reg        [5:0]    io_input_payload_delay_47_partialRound;
  reg        [3:0]    io_input_payload_delay_47_stateIndex;
  reg        [3:0]    io_input_payload_delay_47_stateSize;
  reg        [7:0]    io_input_payload_delay_47_stateID;
  reg        [254:0]  io_input_payload_delay_47_stateElements_0;
  reg        [254:0]  io_input_payload_delay_47_stateElements_1;
  reg        [254:0]  io_input_payload_delay_47_stateElements_2;
  reg        [254:0]  io_input_payload_delay_47_stateElements_3;
  reg        [254:0]  io_input_payload_delay_47_stateElements_4;
  reg        [254:0]  io_input_payload_delay_47_stateElements_5;
  reg        [254:0]  io_input_payload_delay_47_stateElements_6;
  reg        [254:0]  io_input_payload_delay_47_stateElements_7;
  reg        [254:0]  io_input_payload_delay_47_stateElements_8;
  reg        [254:0]  io_input_payload_delay_47_stateElements_9;
  reg        [254:0]  io_input_payload_delay_47_stateElements_10;
  reg        [254:0]  io_input_payload_delay_47_stateElement;
  reg                 io_input_payload_delay_48_isFull;
  reg        [2:0]    io_input_payload_delay_48_fullRound;
  reg        [5:0]    io_input_payload_delay_48_partialRound;
  reg        [3:0]    io_input_payload_delay_48_stateIndex;
  reg        [3:0]    io_input_payload_delay_48_stateSize;
  reg        [7:0]    io_input_payload_delay_48_stateID;
  reg        [254:0]  io_input_payload_delay_48_stateElements_0;
  reg        [254:0]  io_input_payload_delay_48_stateElements_1;
  reg        [254:0]  io_input_payload_delay_48_stateElements_2;
  reg        [254:0]  io_input_payload_delay_48_stateElements_3;
  reg        [254:0]  io_input_payload_delay_48_stateElements_4;
  reg        [254:0]  io_input_payload_delay_48_stateElements_5;
  reg        [254:0]  io_input_payload_delay_48_stateElements_6;
  reg        [254:0]  io_input_payload_delay_48_stateElements_7;
  reg        [254:0]  io_input_payload_delay_48_stateElements_8;
  reg        [254:0]  io_input_payload_delay_48_stateElements_9;
  reg        [254:0]  io_input_payload_delay_48_stateElements_10;
  reg        [254:0]  io_input_payload_delay_48_stateElement;
  reg                 io_input_payload_delay_49_isFull;
  reg        [2:0]    io_input_payload_delay_49_fullRound;
  reg        [5:0]    io_input_payload_delay_49_partialRound;
  reg        [3:0]    io_input_payload_delay_49_stateIndex;
  reg        [3:0]    io_input_payload_delay_49_stateSize;
  reg        [7:0]    io_input_payload_delay_49_stateID;
  reg        [254:0]  io_input_payload_delay_49_stateElements_0;
  reg        [254:0]  io_input_payload_delay_49_stateElements_1;
  reg        [254:0]  io_input_payload_delay_49_stateElements_2;
  reg        [254:0]  io_input_payload_delay_49_stateElements_3;
  reg        [254:0]  io_input_payload_delay_49_stateElements_4;
  reg        [254:0]  io_input_payload_delay_49_stateElements_5;
  reg        [254:0]  io_input_payload_delay_49_stateElements_6;
  reg        [254:0]  io_input_payload_delay_49_stateElements_7;
  reg        [254:0]  io_input_payload_delay_49_stateElements_8;
  reg        [254:0]  io_input_payload_delay_49_stateElements_9;
  reg        [254:0]  io_input_payload_delay_49_stateElements_10;
  reg        [254:0]  io_input_payload_delay_49_stateElement;
  reg                 io_input_payload_delay_50_isFull;
  reg        [2:0]    io_input_payload_delay_50_fullRound;
  reg        [5:0]    io_input_payload_delay_50_partialRound;
  reg        [3:0]    io_input_payload_delay_50_stateIndex;
  reg        [3:0]    io_input_payload_delay_50_stateSize;
  reg        [7:0]    io_input_payload_delay_50_stateID;
  reg        [254:0]  io_input_payload_delay_50_stateElements_0;
  reg        [254:0]  io_input_payload_delay_50_stateElements_1;
  reg        [254:0]  io_input_payload_delay_50_stateElements_2;
  reg        [254:0]  io_input_payload_delay_50_stateElements_3;
  reg        [254:0]  io_input_payload_delay_50_stateElements_4;
  reg        [254:0]  io_input_payload_delay_50_stateElements_5;
  reg        [254:0]  io_input_payload_delay_50_stateElements_6;
  reg        [254:0]  io_input_payload_delay_50_stateElements_7;
  reg        [254:0]  io_input_payload_delay_50_stateElements_8;
  reg        [254:0]  io_input_payload_delay_50_stateElements_9;
  reg        [254:0]  io_input_payload_delay_50_stateElements_10;
  reg        [254:0]  io_input_payload_delay_50_stateElement;
  reg                 io_input_payload_delay_51_isFull;
  reg        [2:0]    io_input_payload_delay_51_fullRound;
  reg        [5:0]    io_input_payload_delay_51_partialRound;
  reg        [3:0]    io_input_payload_delay_51_stateIndex;
  reg        [3:0]    io_input_payload_delay_51_stateSize;
  reg        [7:0]    io_input_payload_delay_51_stateID;
  reg        [254:0]  io_input_payload_delay_51_stateElements_0;
  reg        [254:0]  io_input_payload_delay_51_stateElements_1;
  reg        [254:0]  io_input_payload_delay_51_stateElements_2;
  reg        [254:0]  io_input_payload_delay_51_stateElements_3;
  reg        [254:0]  io_input_payload_delay_51_stateElements_4;
  reg        [254:0]  io_input_payload_delay_51_stateElements_5;
  reg        [254:0]  io_input_payload_delay_51_stateElements_6;
  reg        [254:0]  io_input_payload_delay_51_stateElements_7;
  reg        [254:0]  io_input_payload_delay_51_stateElements_8;
  reg        [254:0]  io_input_payload_delay_51_stateElements_9;
  reg        [254:0]  io_input_payload_delay_51_stateElements_10;
  reg        [254:0]  io_input_payload_delay_51_stateElement;
  reg                 io_input_payload_delay_52_isFull;
  reg        [2:0]    io_input_payload_delay_52_fullRound;
  reg        [5:0]    io_input_payload_delay_52_partialRound;
  reg        [3:0]    io_input_payload_delay_52_stateIndex;
  reg        [3:0]    io_input_payload_delay_52_stateSize;
  reg        [7:0]    io_input_payload_delay_52_stateID;
  reg        [254:0]  io_input_payload_delay_52_stateElements_0;
  reg        [254:0]  io_input_payload_delay_52_stateElements_1;
  reg        [254:0]  io_input_payload_delay_52_stateElements_2;
  reg        [254:0]  io_input_payload_delay_52_stateElements_3;
  reg        [254:0]  io_input_payload_delay_52_stateElements_4;
  reg        [254:0]  io_input_payload_delay_52_stateElements_5;
  reg        [254:0]  io_input_payload_delay_52_stateElements_6;
  reg        [254:0]  io_input_payload_delay_52_stateElements_7;
  reg        [254:0]  io_input_payload_delay_52_stateElements_8;
  reg        [254:0]  io_input_payload_delay_52_stateElements_9;
  reg        [254:0]  io_input_payload_delay_52_stateElements_10;
  reg        [254:0]  io_input_payload_delay_52_stateElement;
  reg                 io_input_payload_delay_53_isFull;
  reg        [2:0]    io_input_payload_delay_53_fullRound;
  reg        [5:0]    io_input_payload_delay_53_partialRound;
  reg        [3:0]    io_input_payload_delay_53_stateIndex;
  reg        [3:0]    io_input_payload_delay_53_stateSize;
  reg        [7:0]    io_input_payload_delay_53_stateID;
  reg        [254:0]  io_input_payload_delay_53_stateElements_0;
  reg        [254:0]  io_input_payload_delay_53_stateElements_1;
  reg        [254:0]  io_input_payload_delay_53_stateElements_2;
  reg        [254:0]  io_input_payload_delay_53_stateElements_3;
  reg        [254:0]  io_input_payload_delay_53_stateElements_4;
  reg        [254:0]  io_input_payload_delay_53_stateElements_5;
  reg        [254:0]  io_input_payload_delay_53_stateElements_6;
  reg        [254:0]  io_input_payload_delay_53_stateElements_7;
  reg        [254:0]  io_input_payload_delay_53_stateElements_8;
  reg        [254:0]  io_input_payload_delay_53_stateElements_9;
  reg        [254:0]  io_input_payload_delay_53_stateElements_10;
  reg        [254:0]  io_input_payload_delay_53_stateElement;
  reg                 io_input_payload_delay_54_isFull;
  reg        [2:0]    io_input_payload_delay_54_fullRound;
  reg        [5:0]    io_input_payload_delay_54_partialRound;
  reg        [3:0]    io_input_payload_delay_54_stateIndex;
  reg        [3:0]    io_input_payload_delay_54_stateSize;
  reg        [7:0]    io_input_payload_delay_54_stateID;
  reg        [254:0]  io_input_payload_delay_54_stateElements_0;
  reg        [254:0]  io_input_payload_delay_54_stateElements_1;
  reg        [254:0]  io_input_payload_delay_54_stateElements_2;
  reg        [254:0]  io_input_payload_delay_54_stateElements_3;
  reg        [254:0]  io_input_payload_delay_54_stateElements_4;
  reg        [254:0]  io_input_payload_delay_54_stateElements_5;
  reg        [254:0]  io_input_payload_delay_54_stateElements_6;
  reg        [254:0]  io_input_payload_delay_54_stateElements_7;
  reg        [254:0]  io_input_payload_delay_54_stateElements_8;
  reg        [254:0]  io_input_payload_delay_54_stateElements_9;
  reg        [254:0]  io_input_payload_delay_54_stateElements_10;
  reg        [254:0]  io_input_payload_delay_54_stateElement;
  reg                 io_input_payload_delay_55_isFull;
  reg        [2:0]    io_input_payload_delay_55_fullRound;
  reg        [5:0]    io_input_payload_delay_55_partialRound;
  reg        [3:0]    io_input_payload_delay_55_stateIndex;
  reg        [3:0]    io_input_payload_delay_55_stateSize;
  reg        [7:0]    io_input_payload_delay_55_stateID;
  reg        [254:0]  io_input_payload_delay_55_stateElements_0;
  reg        [254:0]  io_input_payload_delay_55_stateElements_1;
  reg        [254:0]  io_input_payload_delay_55_stateElements_2;
  reg        [254:0]  io_input_payload_delay_55_stateElements_3;
  reg        [254:0]  io_input_payload_delay_55_stateElements_4;
  reg        [254:0]  io_input_payload_delay_55_stateElements_5;
  reg        [254:0]  io_input_payload_delay_55_stateElements_6;
  reg        [254:0]  io_input_payload_delay_55_stateElements_7;
  reg        [254:0]  io_input_payload_delay_55_stateElements_8;
  reg        [254:0]  io_input_payload_delay_55_stateElements_9;
  reg        [254:0]  io_input_payload_delay_55_stateElements_10;
  reg        [254:0]  io_input_payload_delay_55_stateElement;
  reg                 io_input_payload_delay_56_isFull;
  reg        [2:0]    io_input_payload_delay_56_fullRound;
  reg        [5:0]    io_input_payload_delay_56_partialRound;
  reg        [3:0]    io_input_payload_delay_56_stateIndex;
  reg        [3:0]    io_input_payload_delay_56_stateSize;
  reg        [7:0]    io_input_payload_delay_56_stateID;
  reg        [254:0]  io_input_payload_delay_56_stateElements_0;
  reg        [254:0]  io_input_payload_delay_56_stateElements_1;
  reg        [254:0]  io_input_payload_delay_56_stateElements_2;
  reg        [254:0]  io_input_payload_delay_56_stateElements_3;
  reg        [254:0]  io_input_payload_delay_56_stateElements_4;
  reg        [254:0]  io_input_payload_delay_56_stateElements_5;
  reg        [254:0]  io_input_payload_delay_56_stateElements_6;
  reg        [254:0]  io_input_payload_delay_56_stateElements_7;
  reg        [254:0]  io_input_payload_delay_56_stateElements_8;
  reg        [254:0]  io_input_payload_delay_56_stateElements_9;
  reg        [254:0]  io_input_payload_delay_56_stateElements_10;
  reg        [254:0]  io_input_payload_delay_56_stateElement;
  reg                 io_input_payload_delay_57_isFull;
  reg        [2:0]    io_input_payload_delay_57_fullRound;
  reg        [5:0]    io_input_payload_delay_57_partialRound;
  reg        [3:0]    io_input_payload_delay_57_stateIndex;
  reg        [3:0]    io_input_payload_delay_57_stateSize;
  reg        [7:0]    io_input_payload_delay_57_stateID;
  reg        [254:0]  io_input_payload_delay_57_stateElements_0;
  reg        [254:0]  io_input_payload_delay_57_stateElements_1;
  reg        [254:0]  io_input_payload_delay_57_stateElements_2;
  reg        [254:0]  io_input_payload_delay_57_stateElements_3;
  reg        [254:0]  io_input_payload_delay_57_stateElements_4;
  reg        [254:0]  io_input_payload_delay_57_stateElements_5;
  reg        [254:0]  io_input_payload_delay_57_stateElements_6;
  reg        [254:0]  io_input_payload_delay_57_stateElements_7;
  reg        [254:0]  io_input_payload_delay_57_stateElements_8;
  reg        [254:0]  io_input_payload_delay_57_stateElements_9;
  reg        [254:0]  io_input_payload_delay_57_stateElements_10;
  reg        [254:0]  io_input_payload_delay_57_stateElement;
  reg                 io_input_payload_delay_58_isFull;
  reg        [2:0]    io_input_payload_delay_58_fullRound;
  reg        [5:0]    io_input_payload_delay_58_partialRound;
  reg        [3:0]    io_input_payload_delay_58_stateIndex;
  reg        [3:0]    io_input_payload_delay_58_stateSize;
  reg        [7:0]    io_input_payload_delay_58_stateID;
  reg        [254:0]  io_input_payload_delay_58_stateElements_0;
  reg        [254:0]  io_input_payload_delay_58_stateElements_1;
  reg        [254:0]  io_input_payload_delay_58_stateElements_2;
  reg        [254:0]  io_input_payload_delay_58_stateElements_3;
  reg        [254:0]  io_input_payload_delay_58_stateElements_4;
  reg        [254:0]  io_input_payload_delay_58_stateElements_5;
  reg        [254:0]  io_input_payload_delay_58_stateElements_6;
  reg        [254:0]  io_input_payload_delay_58_stateElements_7;
  reg        [254:0]  io_input_payload_delay_58_stateElements_8;
  reg        [254:0]  io_input_payload_delay_58_stateElements_9;
  reg        [254:0]  io_input_payload_delay_58_stateElements_10;
  reg        [254:0]  io_input_payload_delay_58_stateElement;
  reg                 io_input_payload_delay_59_isFull;
  reg        [2:0]    io_input_payload_delay_59_fullRound;
  reg        [5:0]    io_input_payload_delay_59_partialRound;
  reg        [3:0]    io_input_payload_delay_59_stateIndex;
  reg        [3:0]    io_input_payload_delay_59_stateSize;
  reg        [7:0]    io_input_payload_delay_59_stateID;
  reg        [254:0]  io_input_payload_delay_59_stateElements_0;
  reg        [254:0]  io_input_payload_delay_59_stateElements_1;
  reg        [254:0]  io_input_payload_delay_59_stateElements_2;
  reg        [254:0]  io_input_payload_delay_59_stateElements_3;
  reg        [254:0]  io_input_payload_delay_59_stateElements_4;
  reg        [254:0]  io_input_payload_delay_59_stateElements_5;
  reg        [254:0]  io_input_payload_delay_59_stateElements_6;
  reg        [254:0]  io_input_payload_delay_59_stateElements_7;
  reg        [254:0]  io_input_payload_delay_59_stateElements_8;
  reg        [254:0]  io_input_payload_delay_59_stateElements_9;
  reg        [254:0]  io_input_payload_delay_59_stateElements_10;
  reg        [254:0]  io_input_payload_delay_59_stateElement;
  reg                 io_input_payload_delay_60_isFull;
  reg        [2:0]    io_input_payload_delay_60_fullRound;
  reg        [5:0]    io_input_payload_delay_60_partialRound;
  reg        [3:0]    io_input_payload_delay_60_stateIndex;
  reg        [3:0]    io_input_payload_delay_60_stateSize;
  reg        [7:0]    io_input_payload_delay_60_stateID;
  reg        [254:0]  io_input_payload_delay_60_stateElements_0;
  reg        [254:0]  io_input_payload_delay_60_stateElements_1;
  reg        [254:0]  io_input_payload_delay_60_stateElements_2;
  reg        [254:0]  io_input_payload_delay_60_stateElements_3;
  reg        [254:0]  io_input_payload_delay_60_stateElements_4;
  reg        [254:0]  io_input_payload_delay_60_stateElements_5;
  reg        [254:0]  io_input_payload_delay_60_stateElements_6;
  reg        [254:0]  io_input_payload_delay_60_stateElements_7;
  reg        [254:0]  io_input_payload_delay_60_stateElements_8;
  reg        [254:0]  io_input_payload_delay_60_stateElements_9;
  reg        [254:0]  io_input_payload_delay_60_stateElements_10;
  reg        [254:0]  io_input_payload_delay_60_stateElement;
  reg                 io_input_payload_delay_61_isFull;
  reg        [2:0]    io_input_payload_delay_61_fullRound;
  reg        [5:0]    io_input_payload_delay_61_partialRound;
  reg        [3:0]    io_input_payload_delay_61_stateIndex;
  reg        [3:0]    io_input_payload_delay_61_stateSize;
  reg        [7:0]    io_input_payload_delay_61_stateID;
  reg        [254:0]  io_input_payload_delay_61_stateElements_0;
  reg        [254:0]  io_input_payload_delay_61_stateElements_1;
  reg        [254:0]  io_input_payload_delay_61_stateElements_2;
  reg        [254:0]  io_input_payload_delay_61_stateElements_3;
  reg        [254:0]  io_input_payload_delay_61_stateElements_4;
  reg        [254:0]  io_input_payload_delay_61_stateElements_5;
  reg        [254:0]  io_input_payload_delay_61_stateElements_6;
  reg        [254:0]  io_input_payload_delay_61_stateElements_7;
  reg        [254:0]  io_input_payload_delay_61_stateElements_8;
  reg        [254:0]  io_input_payload_delay_61_stateElements_9;
  reg        [254:0]  io_input_payload_delay_61_stateElements_10;
  reg        [254:0]  io_input_payload_delay_61_stateElement;
  reg                 io_input_payload_delay_62_isFull;
  reg        [2:0]    io_input_payload_delay_62_fullRound;
  reg        [5:0]    io_input_payload_delay_62_partialRound;
  reg        [3:0]    io_input_payload_delay_62_stateIndex;
  reg        [3:0]    io_input_payload_delay_62_stateSize;
  reg        [7:0]    io_input_payload_delay_62_stateID;
  reg        [254:0]  io_input_payload_delay_62_stateElements_0;
  reg        [254:0]  io_input_payload_delay_62_stateElements_1;
  reg        [254:0]  io_input_payload_delay_62_stateElements_2;
  reg        [254:0]  io_input_payload_delay_62_stateElements_3;
  reg        [254:0]  io_input_payload_delay_62_stateElements_4;
  reg        [254:0]  io_input_payload_delay_62_stateElements_5;
  reg        [254:0]  io_input_payload_delay_62_stateElements_6;
  reg        [254:0]  io_input_payload_delay_62_stateElements_7;
  reg        [254:0]  io_input_payload_delay_62_stateElements_8;
  reg        [254:0]  io_input_payload_delay_62_stateElements_9;
  reg        [254:0]  io_input_payload_delay_62_stateElements_10;
  reg        [254:0]  io_input_payload_delay_62_stateElement;
  reg                 io_input_payload_delay_63_isFull;
  reg        [2:0]    io_input_payload_delay_63_fullRound;
  reg        [5:0]    io_input_payload_delay_63_partialRound;
  reg        [3:0]    io_input_payload_delay_63_stateIndex;
  reg        [3:0]    io_input_payload_delay_63_stateSize;
  reg        [7:0]    io_input_payload_delay_63_stateID;
  reg        [254:0]  io_input_payload_delay_63_stateElements_0;
  reg        [254:0]  io_input_payload_delay_63_stateElements_1;
  reg        [254:0]  io_input_payload_delay_63_stateElements_2;
  reg        [254:0]  io_input_payload_delay_63_stateElements_3;
  reg        [254:0]  io_input_payload_delay_63_stateElements_4;
  reg        [254:0]  io_input_payload_delay_63_stateElements_5;
  reg        [254:0]  io_input_payload_delay_63_stateElements_6;
  reg        [254:0]  io_input_payload_delay_63_stateElements_7;
  reg        [254:0]  io_input_payload_delay_63_stateElements_8;
  reg        [254:0]  io_input_payload_delay_63_stateElements_9;
  reg        [254:0]  io_input_payload_delay_63_stateElements_10;
  reg        [254:0]  io_input_payload_delay_63_stateElement;
  reg                 io_input_payload_delay_64_isFull;
  reg        [2:0]    io_input_payload_delay_64_fullRound;
  reg        [5:0]    io_input_payload_delay_64_partialRound;
  reg        [3:0]    io_input_payload_delay_64_stateIndex;
  reg        [3:0]    io_input_payload_delay_64_stateSize;
  reg        [7:0]    io_input_payload_delay_64_stateID;
  reg        [254:0]  io_input_payload_delay_64_stateElements_0;
  reg        [254:0]  io_input_payload_delay_64_stateElements_1;
  reg        [254:0]  io_input_payload_delay_64_stateElements_2;
  reg        [254:0]  io_input_payload_delay_64_stateElements_3;
  reg        [254:0]  io_input_payload_delay_64_stateElements_4;
  reg        [254:0]  io_input_payload_delay_64_stateElements_5;
  reg        [254:0]  io_input_payload_delay_64_stateElements_6;
  reg        [254:0]  io_input_payload_delay_64_stateElements_7;
  reg        [254:0]  io_input_payload_delay_64_stateElements_8;
  reg        [254:0]  io_input_payload_delay_64_stateElements_9;
  reg        [254:0]  io_input_payload_delay_64_stateElements_10;
  reg        [254:0]  io_input_payload_delay_64_stateElement;
  reg                 io_input_payload_delay_65_isFull;
  reg        [2:0]    io_input_payload_delay_65_fullRound;
  reg        [5:0]    io_input_payload_delay_65_partialRound;
  reg        [3:0]    io_input_payload_delay_65_stateIndex;
  reg        [3:0]    io_input_payload_delay_65_stateSize;
  reg        [7:0]    io_input_payload_delay_65_stateID;
  reg        [254:0]  io_input_payload_delay_65_stateElements_0;
  reg        [254:0]  io_input_payload_delay_65_stateElements_1;
  reg        [254:0]  io_input_payload_delay_65_stateElements_2;
  reg        [254:0]  io_input_payload_delay_65_stateElements_3;
  reg        [254:0]  io_input_payload_delay_65_stateElements_4;
  reg        [254:0]  io_input_payload_delay_65_stateElements_5;
  reg        [254:0]  io_input_payload_delay_65_stateElements_6;
  reg        [254:0]  io_input_payload_delay_65_stateElements_7;
  reg        [254:0]  io_input_payload_delay_65_stateElements_8;
  reg        [254:0]  io_input_payload_delay_65_stateElements_9;
  reg        [254:0]  io_input_payload_delay_65_stateElements_10;
  reg        [254:0]  io_input_payload_delay_65_stateElement;
  reg                 io_input_payload_delay_66_isFull;
  reg        [2:0]    io_input_payload_delay_66_fullRound;
  reg        [5:0]    io_input_payload_delay_66_partialRound;
  reg        [3:0]    io_input_payload_delay_66_stateIndex;
  reg        [3:0]    io_input_payload_delay_66_stateSize;
  reg        [7:0]    io_input_payload_delay_66_stateID;
  reg        [254:0]  io_input_payload_delay_66_stateElements_0;
  reg        [254:0]  io_input_payload_delay_66_stateElements_1;
  reg        [254:0]  io_input_payload_delay_66_stateElements_2;
  reg        [254:0]  io_input_payload_delay_66_stateElements_3;
  reg        [254:0]  io_input_payload_delay_66_stateElements_4;
  reg        [254:0]  io_input_payload_delay_66_stateElements_5;
  reg        [254:0]  io_input_payload_delay_66_stateElements_6;
  reg        [254:0]  io_input_payload_delay_66_stateElements_7;
  reg        [254:0]  io_input_payload_delay_66_stateElements_8;
  reg        [254:0]  io_input_payload_delay_66_stateElements_9;
  reg        [254:0]  io_input_payload_delay_66_stateElements_10;
  reg        [254:0]  io_input_payload_delay_66_stateElement;
  reg                 io_input_payload_delay_67_isFull;
  reg        [2:0]    io_input_payload_delay_67_fullRound;
  reg        [5:0]    io_input_payload_delay_67_partialRound;
  reg        [3:0]    io_input_payload_delay_67_stateIndex;
  reg        [3:0]    io_input_payload_delay_67_stateSize;
  reg        [7:0]    io_input_payload_delay_67_stateID;
  reg        [254:0]  io_input_payload_delay_67_stateElements_0;
  reg        [254:0]  io_input_payload_delay_67_stateElements_1;
  reg        [254:0]  io_input_payload_delay_67_stateElements_2;
  reg        [254:0]  io_input_payload_delay_67_stateElements_3;
  reg        [254:0]  io_input_payload_delay_67_stateElements_4;
  reg        [254:0]  io_input_payload_delay_67_stateElements_5;
  reg        [254:0]  io_input_payload_delay_67_stateElements_6;
  reg        [254:0]  io_input_payload_delay_67_stateElements_7;
  reg        [254:0]  io_input_payload_delay_67_stateElements_8;
  reg        [254:0]  io_input_payload_delay_67_stateElements_9;
  reg        [254:0]  io_input_payload_delay_67_stateElements_10;
  reg        [254:0]  io_input_payload_delay_67_stateElement;
  reg                 io_input_payload_delay_68_isFull;
  reg        [2:0]    io_input_payload_delay_68_fullRound;
  reg        [5:0]    io_input_payload_delay_68_partialRound;
  reg        [3:0]    io_input_payload_delay_68_stateIndex;
  reg        [3:0]    io_input_payload_delay_68_stateSize;
  reg        [7:0]    io_input_payload_delay_68_stateID;
  reg        [254:0]  io_input_payload_delay_68_stateElements_0;
  reg        [254:0]  io_input_payload_delay_68_stateElements_1;
  reg        [254:0]  io_input_payload_delay_68_stateElements_2;
  reg        [254:0]  io_input_payload_delay_68_stateElements_3;
  reg        [254:0]  io_input_payload_delay_68_stateElements_4;
  reg        [254:0]  io_input_payload_delay_68_stateElements_5;
  reg        [254:0]  io_input_payload_delay_68_stateElements_6;
  reg        [254:0]  io_input_payload_delay_68_stateElements_7;
  reg        [254:0]  io_input_payload_delay_68_stateElements_8;
  reg        [254:0]  io_input_payload_delay_68_stateElements_9;
  reg        [254:0]  io_input_payload_delay_68_stateElements_10;
  reg        [254:0]  io_input_payload_delay_68_stateElement;
  reg                 io_input_payload_delay_69_isFull;
  reg        [2:0]    io_input_payload_delay_69_fullRound;
  reg        [5:0]    io_input_payload_delay_69_partialRound;
  reg        [3:0]    io_input_payload_delay_69_stateIndex;
  reg        [3:0]    io_input_payload_delay_69_stateSize;
  reg        [7:0]    io_input_payload_delay_69_stateID;
  reg        [254:0]  io_input_payload_delay_69_stateElements_0;
  reg        [254:0]  io_input_payload_delay_69_stateElements_1;
  reg        [254:0]  io_input_payload_delay_69_stateElements_2;
  reg        [254:0]  io_input_payload_delay_69_stateElements_3;
  reg        [254:0]  io_input_payload_delay_69_stateElements_4;
  reg        [254:0]  io_input_payload_delay_69_stateElements_5;
  reg        [254:0]  io_input_payload_delay_69_stateElements_6;
  reg        [254:0]  io_input_payload_delay_69_stateElements_7;
  reg        [254:0]  io_input_payload_delay_69_stateElements_8;
  reg        [254:0]  io_input_payload_delay_69_stateElements_9;
  reg        [254:0]  io_input_payload_delay_69_stateElements_10;
  reg        [254:0]  io_input_payload_delay_69_stateElement;
  reg                 io_input_payload_delay_70_isFull;
  reg        [2:0]    io_input_payload_delay_70_fullRound;
  reg        [5:0]    io_input_payload_delay_70_partialRound;
  reg        [3:0]    io_input_payload_delay_70_stateIndex;
  reg        [3:0]    io_input_payload_delay_70_stateSize;
  reg        [7:0]    io_input_payload_delay_70_stateID;
  reg        [254:0]  io_input_payload_delay_70_stateElements_0;
  reg        [254:0]  io_input_payload_delay_70_stateElements_1;
  reg        [254:0]  io_input_payload_delay_70_stateElements_2;
  reg        [254:0]  io_input_payload_delay_70_stateElements_3;
  reg        [254:0]  io_input_payload_delay_70_stateElements_4;
  reg        [254:0]  io_input_payload_delay_70_stateElements_5;
  reg        [254:0]  io_input_payload_delay_70_stateElements_6;
  reg        [254:0]  io_input_payload_delay_70_stateElements_7;
  reg        [254:0]  io_input_payload_delay_70_stateElements_8;
  reg        [254:0]  io_input_payload_delay_70_stateElements_9;
  reg        [254:0]  io_input_payload_delay_70_stateElements_10;
  reg        [254:0]  io_input_payload_delay_70_stateElement;
  reg                 io_input_payload_delay_71_isFull;
  reg        [2:0]    io_input_payload_delay_71_fullRound;
  reg        [5:0]    io_input_payload_delay_71_partialRound;
  reg        [3:0]    io_input_payload_delay_71_stateIndex;
  reg        [3:0]    io_input_payload_delay_71_stateSize;
  reg        [7:0]    io_input_payload_delay_71_stateID;
  reg        [254:0]  io_input_payload_delay_71_stateElements_0;
  reg        [254:0]  io_input_payload_delay_71_stateElements_1;
  reg        [254:0]  io_input_payload_delay_71_stateElements_2;
  reg        [254:0]  io_input_payload_delay_71_stateElements_3;
  reg        [254:0]  io_input_payload_delay_71_stateElements_4;
  reg        [254:0]  io_input_payload_delay_71_stateElements_5;
  reg        [254:0]  io_input_payload_delay_71_stateElements_6;
  reg        [254:0]  io_input_payload_delay_71_stateElements_7;
  reg        [254:0]  io_input_payload_delay_71_stateElements_8;
  reg        [254:0]  io_input_payload_delay_71_stateElements_9;
  reg        [254:0]  io_input_payload_delay_71_stateElements_10;
  reg        [254:0]  io_input_payload_delay_71_stateElement;
  reg                 io_input_payload_delay_72_isFull;
  reg        [2:0]    io_input_payload_delay_72_fullRound;
  reg        [5:0]    io_input_payload_delay_72_partialRound;
  reg        [3:0]    io_input_payload_delay_72_stateIndex;
  reg        [3:0]    io_input_payload_delay_72_stateSize;
  reg        [7:0]    io_input_payload_delay_72_stateID;
  reg        [254:0]  io_input_payload_delay_72_stateElements_0;
  reg        [254:0]  io_input_payload_delay_72_stateElements_1;
  reg        [254:0]  io_input_payload_delay_72_stateElements_2;
  reg        [254:0]  io_input_payload_delay_72_stateElements_3;
  reg        [254:0]  io_input_payload_delay_72_stateElements_4;
  reg        [254:0]  io_input_payload_delay_72_stateElements_5;
  reg        [254:0]  io_input_payload_delay_72_stateElements_6;
  reg        [254:0]  io_input_payload_delay_72_stateElements_7;
  reg        [254:0]  io_input_payload_delay_72_stateElements_8;
  reg        [254:0]  io_input_payload_delay_72_stateElements_9;
  reg        [254:0]  io_input_payload_delay_72_stateElements_10;
  reg        [254:0]  io_input_payload_delay_72_stateElement;
  reg                 io_input_payload_delay_73_isFull;
  reg        [2:0]    io_input_payload_delay_73_fullRound;
  reg        [5:0]    io_input_payload_delay_73_partialRound;
  reg        [3:0]    io_input_payload_delay_73_stateIndex;
  reg        [3:0]    io_input_payload_delay_73_stateSize;
  reg        [7:0]    io_input_payload_delay_73_stateID;
  reg        [254:0]  io_input_payload_delay_73_stateElements_0;
  reg        [254:0]  io_input_payload_delay_73_stateElements_1;
  reg        [254:0]  io_input_payload_delay_73_stateElements_2;
  reg        [254:0]  io_input_payload_delay_73_stateElements_3;
  reg        [254:0]  io_input_payload_delay_73_stateElements_4;
  reg        [254:0]  io_input_payload_delay_73_stateElements_5;
  reg        [254:0]  io_input_payload_delay_73_stateElements_6;
  reg        [254:0]  io_input_payload_delay_73_stateElements_7;
  reg        [254:0]  io_input_payload_delay_73_stateElements_8;
  reg        [254:0]  io_input_payload_delay_73_stateElements_9;
  reg        [254:0]  io_input_payload_delay_73_stateElements_10;
  reg        [254:0]  io_input_payload_delay_73_stateElement;
  reg                 io_input_payload_delay_74_isFull;
  reg        [2:0]    io_input_payload_delay_74_fullRound;
  reg        [5:0]    io_input_payload_delay_74_partialRound;
  reg        [3:0]    io_input_payload_delay_74_stateIndex;
  reg        [3:0]    io_input_payload_delay_74_stateSize;
  reg        [7:0]    io_input_payload_delay_74_stateID;
  reg        [254:0]  io_input_payload_delay_74_stateElements_0;
  reg        [254:0]  io_input_payload_delay_74_stateElements_1;
  reg        [254:0]  io_input_payload_delay_74_stateElements_2;
  reg        [254:0]  io_input_payload_delay_74_stateElements_3;
  reg        [254:0]  io_input_payload_delay_74_stateElements_4;
  reg        [254:0]  io_input_payload_delay_74_stateElements_5;
  reg        [254:0]  io_input_payload_delay_74_stateElements_6;
  reg        [254:0]  io_input_payload_delay_74_stateElements_7;
  reg        [254:0]  io_input_payload_delay_74_stateElements_8;
  reg        [254:0]  io_input_payload_delay_74_stateElements_9;
  reg        [254:0]  io_input_payload_delay_74_stateElements_10;
  reg        [254:0]  io_input_payload_delay_74_stateElement;
  reg                 io_input_payload_delay_75_isFull;
  reg        [2:0]    io_input_payload_delay_75_fullRound;
  reg        [5:0]    io_input_payload_delay_75_partialRound;
  reg        [3:0]    io_input_payload_delay_75_stateIndex;
  reg        [3:0]    io_input_payload_delay_75_stateSize;
  reg        [7:0]    io_input_payload_delay_75_stateID;
  reg        [254:0]  io_input_payload_delay_75_stateElements_0;
  reg        [254:0]  io_input_payload_delay_75_stateElements_1;
  reg        [254:0]  io_input_payload_delay_75_stateElements_2;
  reg        [254:0]  io_input_payload_delay_75_stateElements_3;
  reg        [254:0]  io_input_payload_delay_75_stateElements_4;
  reg        [254:0]  io_input_payload_delay_75_stateElements_5;
  reg        [254:0]  io_input_payload_delay_75_stateElements_6;
  reg        [254:0]  io_input_payload_delay_75_stateElements_7;
  reg        [254:0]  io_input_payload_delay_75_stateElements_8;
  reg        [254:0]  io_input_payload_delay_75_stateElements_9;
  reg        [254:0]  io_input_payload_delay_75_stateElements_10;
  reg        [254:0]  io_input_payload_delay_75_stateElement;
  reg                 io_input_payload_delay_76_isFull;
  reg        [2:0]    io_input_payload_delay_76_fullRound;
  reg        [5:0]    io_input_payload_delay_76_partialRound;
  reg        [3:0]    io_input_payload_delay_76_stateIndex;
  reg        [3:0]    io_input_payload_delay_76_stateSize;
  reg        [7:0]    io_input_payload_delay_76_stateID;
  reg        [254:0]  io_input_payload_delay_76_stateElements_0;
  reg        [254:0]  io_input_payload_delay_76_stateElements_1;
  reg        [254:0]  io_input_payload_delay_76_stateElements_2;
  reg        [254:0]  io_input_payload_delay_76_stateElements_3;
  reg        [254:0]  io_input_payload_delay_76_stateElements_4;
  reg        [254:0]  io_input_payload_delay_76_stateElements_5;
  reg        [254:0]  io_input_payload_delay_76_stateElements_6;
  reg        [254:0]  io_input_payload_delay_76_stateElements_7;
  reg        [254:0]  io_input_payload_delay_76_stateElements_8;
  reg        [254:0]  io_input_payload_delay_76_stateElements_9;
  reg        [254:0]  io_input_payload_delay_76_stateElements_10;
  reg        [254:0]  io_input_payload_delay_76_stateElement;
  reg                 io_input_payload_delay_77_isFull;
  reg        [2:0]    io_input_payload_delay_77_fullRound;
  reg        [5:0]    io_input_payload_delay_77_partialRound;
  reg        [3:0]    io_input_payload_delay_77_stateIndex;
  reg        [3:0]    io_input_payload_delay_77_stateSize;
  reg        [7:0]    io_input_payload_delay_77_stateID;
  reg        [254:0]  io_input_payload_delay_77_stateElements_0;
  reg        [254:0]  io_input_payload_delay_77_stateElements_1;
  reg        [254:0]  io_input_payload_delay_77_stateElements_2;
  reg        [254:0]  io_input_payload_delay_77_stateElements_3;
  reg        [254:0]  io_input_payload_delay_77_stateElements_4;
  reg        [254:0]  io_input_payload_delay_77_stateElements_5;
  reg        [254:0]  io_input_payload_delay_77_stateElements_6;
  reg        [254:0]  io_input_payload_delay_77_stateElements_7;
  reg        [254:0]  io_input_payload_delay_77_stateElements_8;
  reg        [254:0]  io_input_payload_delay_77_stateElements_9;
  reg        [254:0]  io_input_payload_delay_77_stateElements_10;
  reg        [254:0]  io_input_payload_delay_77_stateElement;
  reg                 io_input_payload_delay_78_isFull;
  reg        [2:0]    io_input_payload_delay_78_fullRound;
  reg        [5:0]    io_input_payload_delay_78_partialRound;
  reg        [3:0]    io_input_payload_delay_78_stateIndex;
  reg        [3:0]    io_input_payload_delay_78_stateSize;
  reg        [7:0]    io_input_payload_delay_78_stateID;
  reg        [254:0]  io_input_payload_delay_78_stateElements_0;
  reg        [254:0]  io_input_payload_delay_78_stateElements_1;
  reg        [254:0]  io_input_payload_delay_78_stateElements_2;
  reg        [254:0]  io_input_payload_delay_78_stateElements_3;
  reg        [254:0]  io_input_payload_delay_78_stateElements_4;
  reg        [254:0]  io_input_payload_delay_78_stateElements_5;
  reg        [254:0]  io_input_payload_delay_78_stateElements_6;
  reg        [254:0]  io_input_payload_delay_78_stateElements_7;
  reg        [254:0]  io_input_payload_delay_78_stateElements_8;
  reg        [254:0]  io_input_payload_delay_78_stateElements_9;
  reg        [254:0]  io_input_payload_delay_78_stateElements_10;
  reg        [254:0]  io_input_payload_delay_78_stateElement;
  reg                 io_input_payload_delay_79_isFull;
  reg        [2:0]    io_input_payload_delay_79_fullRound;
  reg        [5:0]    io_input_payload_delay_79_partialRound;
  reg        [3:0]    io_input_payload_delay_79_stateIndex;
  reg        [3:0]    io_input_payload_delay_79_stateSize;
  reg        [7:0]    io_input_payload_delay_79_stateID;
  reg        [254:0]  io_input_payload_delay_79_stateElements_0;
  reg        [254:0]  io_input_payload_delay_79_stateElements_1;
  reg        [254:0]  io_input_payload_delay_79_stateElements_2;
  reg        [254:0]  io_input_payload_delay_79_stateElements_3;
  reg        [254:0]  io_input_payload_delay_79_stateElements_4;
  reg        [254:0]  io_input_payload_delay_79_stateElements_5;
  reg        [254:0]  io_input_payload_delay_79_stateElements_6;
  reg        [254:0]  io_input_payload_delay_79_stateElements_7;
  reg        [254:0]  io_input_payload_delay_79_stateElements_8;
  reg        [254:0]  io_input_payload_delay_79_stateElements_9;
  reg        [254:0]  io_input_payload_delay_79_stateElements_10;
  reg        [254:0]  io_input_payload_delay_79_stateElement;
  reg                 io_input_payload_delay_80_isFull;
  reg        [2:0]    io_input_payload_delay_80_fullRound;
  reg        [5:0]    io_input_payload_delay_80_partialRound;
  reg        [3:0]    io_input_payload_delay_80_stateIndex;
  reg        [3:0]    io_input_payload_delay_80_stateSize;
  reg        [7:0]    io_input_payload_delay_80_stateID;
  reg        [254:0]  io_input_payload_delay_80_stateElements_0;
  reg        [254:0]  io_input_payload_delay_80_stateElements_1;
  reg        [254:0]  io_input_payload_delay_80_stateElements_2;
  reg        [254:0]  io_input_payload_delay_80_stateElements_3;
  reg        [254:0]  io_input_payload_delay_80_stateElements_4;
  reg        [254:0]  io_input_payload_delay_80_stateElements_5;
  reg        [254:0]  io_input_payload_delay_80_stateElements_6;
  reg        [254:0]  io_input_payload_delay_80_stateElements_7;
  reg        [254:0]  io_input_payload_delay_80_stateElements_8;
  reg        [254:0]  io_input_payload_delay_80_stateElements_9;
  reg        [254:0]  io_input_payload_delay_80_stateElements_10;
  reg        [254:0]  io_input_payload_delay_80_stateElement;
  reg                 io_input_payload_delay_81_isFull;
  reg        [2:0]    io_input_payload_delay_81_fullRound;
  reg        [5:0]    io_input_payload_delay_81_partialRound;
  reg        [3:0]    io_input_payload_delay_81_stateIndex;
  reg        [3:0]    io_input_payload_delay_81_stateSize;
  reg        [7:0]    io_input_payload_delay_81_stateID;
  reg        [254:0]  io_input_payload_delay_81_stateElements_0;
  reg        [254:0]  io_input_payload_delay_81_stateElements_1;
  reg        [254:0]  io_input_payload_delay_81_stateElements_2;
  reg        [254:0]  io_input_payload_delay_81_stateElements_3;
  reg        [254:0]  io_input_payload_delay_81_stateElements_4;
  reg        [254:0]  io_input_payload_delay_81_stateElements_5;
  reg        [254:0]  io_input_payload_delay_81_stateElements_6;
  reg        [254:0]  io_input_payload_delay_81_stateElements_7;
  reg        [254:0]  io_input_payload_delay_81_stateElements_8;
  reg        [254:0]  io_input_payload_delay_81_stateElements_9;
  reg        [254:0]  io_input_payload_delay_81_stateElements_10;
  reg        [254:0]  io_input_payload_delay_81_stateElement;
  reg                 io_input_payload_delay_82_isFull;
  reg        [2:0]    io_input_payload_delay_82_fullRound;
  reg        [5:0]    io_input_payload_delay_82_partialRound;
  reg        [3:0]    io_input_payload_delay_82_stateIndex;
  reg        [3:0]    io_input_payload_delay_82_stateSize;
  reg        [7:0]    io_input_payload_delay_82_stateID;
  reg        [254:0]  io_input_payload_delay_82_stateElements_0;
  reg        [254:0]  io_input_payload_delay_82_stateElements_1;
  reg        [254:0]  io_input_payload_delay_82_stateElements_2;
  reg        [254:0]  io_input_payload_delay_82_stateElements_3;
  reg        [254:0]  io_input_payload_delay_82_stateElements_4;
  reg        [254:0]  io_input_payload_delay_82_stateElements_5;
  reg        [254:0]  io_input_payload_delay_82_stateElements_6;
  reg        [254:0]  io_input_payload_delay_82_stateElements_7;
  reg        [254:0]  io_input_payload_delay_82_stateElements_8;
  reg        [254:0]  io_input_payload_delay_82_stateElements_9;
  reg        [254:0]  io_input_payload_delay_82_stateElements_10;
  reg        [254:0]  io_input_payload_delay_82_stateElement;
  reg                 io_input_payload_delay_83_isFull;
  reg        [2:0]    io_input_payload_delay_83_fullRound;
  reg        [5:0]    io_input_payload_delay_83_partialRound;
  reg        [3:0]    io_input_payload_delay_83_stateIndex;
  reg        [3:0]    io_input_payload_delay_83_stateSize;
  reg        [7:0]    io_input_payload_delay_83_stateID;
  reg        [254:0]  io_input_payload_delay_83_stateElements_0;
  reg        [254:0]  io_input_payload_delay_83_stateElements_1;
  reg        [254:0]  io_input_payload_delay_83_stateElements_2;
  reg        [254:0]  io_input_payload_delay_83_stateElements_3;
  reg        [254:0]  io_input_payload_delay_83_stateElements_4;
  reg        [254:0]  io_input_payload_delay_83_stateElements_5;
  reg        [254:0]  io_input_payload_delay_83_stateElements_6;
  reg        [254:0]  io_input_payload_delay_83_stateElements_7;
  reg        [254:0]  io_input_payload_delay_83_stateElements_8;
  reg        [254:0]  io_input_payload_delay_83_stateElements_9;
  reg        [254:0]  io_input_payload_delay_83_stateElements_10;
  reg        [254:0]  io_input_payload_delay_83_stateElement;
  reg                 io_input_payload_delay_84_isFull;
  reg        [2:0]    io_input_payload_delay_84_fullRound;
  reg        [5:0]    io_input_payload_delay_84_partialRound;
  reg        [3:0]    io_input_payload_delay_84_stateIndex;
  reg        [3:0]    io_input_payload_delay_84_stateSize;
  reg        [7:0]    io_input_payload_delay_84_stateID;
  reg        [254:0]  io_input_payload_delay_84_stateElements_0;
  reg        [254:0]  io_input_payload_delay_84_stateElements_1;
  reg        [254:0]  io_input_payload_delay_84_stateElements_2;
  reg        [254:0]  io_input_payload_delay_84_stateElements_3;
  reg        [254:0]  io_input_payload_delay_84_stateElements_4;
  reg        [254:0]  io_input_payload_delay_84_stateElements_5;
  reg        [254:0]  io_input_payload_delay_84_stateElements_6;
  reg        [254:0]  io_input_payload_delay_84_stateElements_7;
  reg        [254:0]  io_input_payload_delay_84_stateElements_8;
  reg        [254:0]  io_input_payload_delay_84_stateElements_9;
  reg        [254:0]  io_input_payload_delay_84_stateElements_10;
  reg        [254:0]  io_input_payload_delay_84_stateElement;
  reg                 io_input_payload_delay_85_isFull;
  reg        [2:0]    io_input_payload_delay_85_fullRound;
  reg        [5:0]    io_input_payload_delay_85_partialRound;
  reg        [3:0]    io_input_payload_delay_85_stateIndex;
  reg        [3:0]    io_input_payload_delay_85_stateSize;
  reg        [7:0]    io_input_payload_delay_85_stateID;
  reg        [254:0]  io_input_payload_delay_85_stateElements_0;
  reg        [254:0]  io_input_payload_delay_85_stateElements_1;
  reg        [254:0]  io_input_payload_delay_85_stateElements_2;
  reg        [254:0]  io_input_payload_delay_85_stateElements_3;
  reg        [254:0]  io_input_payload_delay_85_stateElements_4;
  reg        [254:0]  io_input_payload_delay_85_stateElements_5;
  reg        [254:0]  io_input_payload_delay_85_stateElements_6;
  reg        [254:0]  io_input_payload_delay_85_stateElements_7;
  reg        [254:0]  io_input_payload_delay_85_stateElements_8;
  reg        [254:0]  io_input_payload_delay_85_stateElements_9;
  reg        [254:0]  io_input_payload_delay_85_stateElements_10;
  reg        [254:0]  io_input_payload_delay_85_stateElement;
  reg                 io_input_payload_delay_86_isFull;
  reg        [2:0]    io_input_payload_delay_86_fullRound;
  reg        [5:0]    io_input_payload_delay_86_partialRound;
  reg        [3:0]    io_input_payload_delay_86_stateIndex;
  reg        [3:0]    io_input_payload_delay_86_stateSize;
  reg        [7:0]    io_input_payload_delay_86_stateID;
  reg        [254:0]  io_input_payload_delay_86_stateElements_0;
  reg        [254:0]  io_input_payload_delay_86_stateElements_1;
  reg        [254:0]  io_input_payload_delay_86_stateElements_2;
  reg        [254:0]  io_input_payload_delay_86_stateElements_3;
  reg        [254:0]  io_input_payload_delay_86_stateElements_4;
  reg        [254:0]  io_input_payload_delay_86_stateElements_5;
  reg        [254:0]  io_input_payload_delay_86_stateElements_6;
  reg        [254:0]  io_input_payload_delay_86_stateElements_7;
  reg        [254:0]  io_input_payload_delay_86_stateElements_8;
  reg        [254:0]  io_input_payload_delay_86_stateElements_9;
  reg        [254:0]  io_input_payload_delay_86_stateElements_10;
  reg        [254:0]  io_input_payload_delay_86_stateElement;
  reg                 io_input_payload_delay_87_isFull;
  reg        [2:0]    io_input_payload_delay_87_fullRound;
  reg        [5:0]    io_input_payload_delay_87_partialRound;
  reg        [3:0]    io_input_payload_delay_87_stateIndex;
  reg        [3:0]    io_input_payload_delay_87_stateSize;
  reg        [7:0]    io_input_payload_delay_87_stateID;
  reg        [254:0]  io_input_payload_delay_87_stateElements_0;
  reg        [254:0]  io_input_payload_delay_87_stateElements_1;
  reg        [254:0]  io_input_payload_delay_87_stateElements_2;
  reg        [254:0]  io_input_payload_delay_87_stateElements_3;
  reg        [254:0]  io_input_payload_delay_87_stateElements_4;
  reg        [254:0]  io_input_payload_delay_87_stateElements_5;
  reg        [254:0]  io_input_payload_delay_87_stateElements_6;
  reg        [254:0]  io_input_payload_delay_87_stateElements_7;
  reg        [254:0]  io_input_payload_delay_87_stateElements_8;
  reg        [254:0]  io_input_payload_delay_87_stateElements_9;
  reg        [254:0]  io_input_payload_delay_87_stateElements_10;
  reg        [254:0]  io_input_payload_delay_87_stateElement;
  reg                 io_input_payload_delay_88_isFull;
  reg        [2:0]    io_input_payload_delay_88_fullRound;
  reg        [5:0]    io_input_payload_delay_88_partialRound;
  reg        [3:0]    io_input_payload_delay_88_stateIndex;
  reg        [3:0]    io_input_payload_delay_88_stateSize;
  reg        [7:0]    io_input_payload_delay_88_stateID;
  reg        [254:0]  io_input_payload_delay_88_stateElements_0;
  reg        [254:0]  io_input_payload_delay_88_stateElements_1;
  reg        [254:0]  io_input_payload_delay_88_stateElements_2;
  reg        [254:0]  io_input_payload_delay_88_stateElements_3;
  reg        [254:0]  io_input_payload_delay_88_stateElements_4;
  reg        [254:0]  io_input_payload_delay_88_stateElements_5;
  reg        [254:0]  io_input_payload_delay_88_stateElements_6;
  reg        [254:0]  io_input_payload_delay_88_stateElements_7;
  reg        [254:0]  io_input_payload_delay_88_stateElements_8;
  reg        [254:0]  io_input_payload_delay_88_stateElements_9;
  reg        [254:0]  io_input_payload_delay_88_stateElements_10;
  reg        [254:0]  io_input_payload_delay_88_stateElement;
  reg                 io_input_payload_delay_89_isFull;
  reg        [2:0]    io_input_payload_delay_89_fullRound;
  reg        [5:0]    io_input_payload_delay_89_partialRound;
  reg        [3:0]    io_input_payload_delay_89_stateIndex;
  reg        [3:0]    io_input_payload_delay_89_stateSize;
  reg        [7:0]    io_input_payload_delay_89_stateID;
  reg        [254:0]  io_input_payload_delay_89_stateElements_0;
  reg        [254:0]  io_input_payload_delay_89_stateElements_1;
  reg        [254:0]  io_input_payload_delay_89_stateElements_2;
  reg        [254:0]  io_input_payload_delay_89_stateElements_3;
  reg        [254:0]  io_input_payload_delay_89_stateElements_4;
  reg        [254:0]  io_input_payload_delay_89_stateElements_5;
  reg        [254:0]  io_input_payload_delay_89_stateElements_6;
  reg        [254:0]  io_input_payload_delay_89_stateElements_7;
  reg        [254:0]  io_input_payload_delay_89_stateElements_8;
  reg        [254:0]  io_input_payload_delay_89_stateElements_9;
  reg        [254:0]  io_input_payload_delay_89_stateElements_10;
  reg        [254:0]  io_input_payload_delay_89_stateElement;
  reg                 io_input_payload_delay_90_isFull;
  reg        [2:0]    io_input_payload_delay_90_fullRound;
  reg        [5:0]    io_input_payload_delay_90_partialRound;
  reg        [3:0]    io_input_payload_delay_90_stateIndex;
  reg        [3:0]    io_input_payload_delay_90_stateSize;
  reg        [7:0]    io_input_payload_delay_90_stateID;
  reg        [254:0]  io_input_payload_delay_90_stateElements_0;
  reg        [254:0]  io_input_payload_delay_90_stateElements_1;
  reg        [254:0]  io_input_payload_delay_90_stateElements_2;
  reg        [254:0]  io_input_payload_delay_90_stateElements_3;
  reg        [254:0]  io_input_payload_delay_90_stateElements_4;
  reg        [254:0]  io_input_payload_delay_90_stateElements_5;
  reg        [254:0]  io_input_payload_delay_90_stateElements_6;
  reg        [254:0]  io_input_payload_delay_90_stateElements_7;
  reg        [254:0]  io_input_payload_delay_90_stateElements_8;
  reg        [254:0]  io_input_payload_delay_90_stateElements_9;
  reg        [254:0]  io_input_payload_delay_90_stateElements_10;
  reg        [254:0]  io_input_payload_delay_90_stateElement;
  reg                 io_input_payload_delay_91_isFull;
  reg        [2:0]    io_input_payload_delay_91_fullRound;
  reg        [5:0]    io_input_payload_delay_91_partialRound;
  reg        [3:0]    io_input_payload_delay_91_stateIndex;
  reg        [3:0]    io_input_payload_delay_91_stateSize;
  reg        [7:0]    io_input_payload_delay_91_stateID;
  reg        [254:0]  io_input_payload_delay_91_stateElements_0;
  reg        [254:0]  io_input_payload_delay_91_stateElements_1;
  reg        [254:0]  io_input_payload_delay_91_stateElements_2;
  reg        [254:0]  io_input_payload_delay_91_stateElements_3;
  reg        [254:0]  io_input_payload_delay_91_stateElements_4;
  reg        [254:0]  io_input_payload_delay_91_stateElements_5;
  reg        [254:0]  io_input_payload_delay_91_stateElements_6;
  reg        [254:0]  io_input_payload_delay_91_stateElements_7;
  reg        [254:0]  io_input_payload_delay_91_stateElements_8;
  reg        [254:0]  io_input_payload_delay_91_stateElements_9;
  reg        [254:0]  io_input_payload_delay_91_stateElements_10;
  reg        [254:0]  io_input_payload_delay_91_stateElement;
  reg                 io_input_payload_delay_92_isFull;
  reg        [2:0]    io_input_payload_delay_92_fullRound;
  reg        [5:0]    io_input_payload_delay_92_partialRound;
  reg        [3:0]    io_input_payload_delay_92_stateIndex;
  reg        [3:0]    io_input_payload_delay_92_stateSize;
  reg        [7:0]    io_input_payload_delay_92_stateID;
  reg        [254:0]  io_input_payload_delay_92_stateElements_0;
  reg        [254:0]  io_input_payload_delay_92_stateElements_1;
  reg        [254:0]  io_input_payload_delay_92_stateElements_2;
  reg        [254:0]  io_input_payload_delay_92_stateElements_3;
  reg        [254:0]  io_input_payload_delay_92_stateElements_4;
  reg        [254:0]  io_input_payload_delay_92_stateElements_5;
  reg        [254:0]  io_input_payload_delay_92_stateElements_6;
  reg        [254:0]  io_input_payload_delay_92_stateElements_7;
  reg        [254:0]  io_input_payload_delay_92_stateElements_8;
  reg        [254:0]  io_input_payload_delay_92_stateElements_9;
  reg        [254:0]  io_input_payload_delay_92_stateElements_10;
  reg        [254:0]  io_input_payload_delay_92_stateElement;
  reg                 io_input_payload_delay_93_isFull;
  reg        [2:0]    io_input_payload_delay_93_fullRound;
  reg        [5:0]    io_input_payload_delay_93_partialRound;
  reg        [3:0]    io_input_payload_delay_93_stateIndex;
  reg        [3:0]    io_input_payload_delay_93_stateSize;
  reg        [7:0]    io_input_payload_delay_93_stateID;
  reg        [254:0]  io_input_payload_delay_93_stateElements_0;
  reg        [254:0]  io_input_payload_delay_93_stateElements_1;
  reg        [254:0]  io_input_payload_delay_93_stateElements_2;
  reg        [254:0]  io_input_payload_delay_93_stateElements_3;
  reg        [254:0]  io_input_payload_delay_93_stateElements_4;
  reg        [254:0]  io_input_payload_delay_93_stateElements_5;
  reg        [254:0]  io_input_payload_delay_93_stateElements_6;
  reg        [254:0]  io_input_payload_delay_93_stateElements_7;
  reg        [254:0]  io_input_payload_delay_93_stateElements_8;
  reg        [254:0]  io_input_payload_delay_93_stateElements_9;
  reg        [254:0]  io_input_payload_delay_93_stateElements_10;
  reg        [254:0]  io_input_payload_delay_93_stateElement;
  reg                 io_input_payload_delay_94_isFull;
  reg        [2:0]    io_input_payload_delay_94_fullRound;
  reg        [5:0]    io_input_payload_delay_94_partialRound;
  reg        [3:0]    io_input_payload_delay_94_stateIndex;
  reg        [3:0]    io_input_payload_delay_94_stateSize;
  reg        [7:0]    io_input_payload_delay_94_stateID;
  reg        [254:0]  io_input_payload_delay_94_stateElements_0;
  reg        [254:0]  io_input_payload_delay_94_stateElements_1;
  reg        [254:0]  io_input_payload_delay_94_stateElements_2;
  reg        [254:0]  io_input_payload_delay_94_stateElements_3;
  reg        [254:0]  io_input_payload_delay_94_stateElements_4;
  reg        [254:0]  io_input_payload_delay_94_stateElements_5;
  reg        [254:0]  io_input_payload_delay_94_stateElements_6;
  reg        [254:0]  io_input_payload_delay_94_stateElements_7;
  reg        [254:0]  io_input_payload_delay_94_stateElements_8;
  reg        [254:0]  io_input_payload_delay_94_stateElements_9;
  reg        [254:0]  io_input_payload_delay_94_stateElements_10;
  reg        [254:0]  io_input_payload_delay_94_stateElement;
  reg                 io_input_payload_delay_95_isFull;
  reg        [2:0]    io_input_payload_delay_95_fullRound;
  reg        [5:0]    io_input_payload_delay_95_partialRound;
  reg        [3:0]    io_input_payload_delay_95_stateIndex;
  reg        [3:0]    io_input_payload_delay_95_stateSize;
  reg        [7:0]    io_input_payload_delay_95_stateID;
  reg        [254:0]  io_input_payload_delay_95_stateElements_0;
  reg        [254:0]  io_input_payload_delay_95_stateElements_1;
  reg        [254:0]  io_input_payload_delay_95_stateElements_2;
  reg        [254:0]  io_input_payload_delay_95_stateElements_3;
  reg        [254:0]  io_input_payload_delay_95_stateElements_4;
  reg        [254:0]  io_input_payload_delay_95_stateElements_5;
  reg        [254:0]  io_input_payload_delay_95_stateElements_6;
  reg        [254:0]  io_input_payload_delay_95_stateElements_7;
  reg        [254:0]  io_input_payload_delay_95_stateElements_8;
  reg        [254:0]  io_input_payload_delay_95_stateElements_9;
  reg        [254:0]  io_input_payload_delay_95_stateElements_10;
  reg        [254:0]  io_input_payload_delay_95_stateElement;
  reg                 io_input_payload_delay_96_isFull;
  reg        [2:0]    io_input_payload_delay_96_fullRound;
  reg        [5:0]    io_input_payload_delay_96_partialRound;
  reg        [3:0]    io_input_payload_delay_96_stateIndex;
  reg        [3:0]    io_input_payload_delay_96_stateSize;
  reg        [7:0]    io_input_payload_delay_96_stateID;
  reg        [254:0]  io_input_payload_delay_96_stateElements_0;
  reg        [254:0]  io_input_payload_delay_96_stateElements_1;
  reg        [254:0]  io_input_payload_delay_96_stateElements_2;
  reg        [254:0]  io_input_payload_delay_96_stateElements_3;
  reg        [254:0]  io_input_payload_delay_96_stateElements_4;
  reg        [254:0]  io_input_payload_delay_96_stateElements_5;
  reg        [254:0]  io_input_payload_delay_96_stateElements_6;
  reg        [254:0]  io_input_payload_delay_96_stateElements_7;
  reg        [254:0]  io_input_payload_delay_96_stateElements_8;
  reg        [254:0]  io_input_payload_delay_96_stateElements_9;
  reg        [254:0]  io_input_payload_delay_96_stateElements_10;
  reg        [254:0]  io_input_payload_delay_96_stateElement;
  reg                 io_input_payload_delay_97_isFull;
  reg        [2:0]    io_input_payload_delay_97_fullRound;
  reg        [5:0]    io_input_payload_delay_97_partialRound;
  reg        [3:0]    io_input_payload_delay_97_stateIndex;
  reg        [3:0]    io_input_payload_delay_97_stateSize;
  reg        [7:0]    io_input_payload_delay_97_stateID;
  reg        [254:0]  io_input_payload_delay_97_stateElements_0;
  reg        [254:0]  io_input_payload_delay_97_stateElements_1;
  reg        [254:0]  io_input_payload_delay_97_stateElements_2;
  reg        [254:0]  io_input_payload_delay_97_stateElements_3;
  reg        [254:0]  io_input_payload_delay_97_stateElements_4;
  reg        [254:0]  io_input_payload_delay_97_stateElements_5;
  reg        [254:0]  io_input_payload_delay_97_stateElements_6;
  reg        [254:0]  io_input_payload_delay_97_stateElements_7;
  reg        [254:0]  io_input_payload_delay_97_stateElements_8;
  reg        [254:0]  io_input_payload_delay_97_stateElements_9;
  reg        [254:0]  io_input_payload_delay_97_stateElements_10;
  reg        [254:0]  io_input_payload_delay_97_stateElement;
  reg                 SBox5Stage_tempContext1_isFull;
  reg        [2:0]    SBox5Stage_tempContext1_fullRound;
  reg        [5:0]    SBox5Stage_tempContext1_partialRound;
  reg        [3:0]    SBox5Stage_tempContext1_stateIndex;
  reg        [3:0]    SBox5Stage_tempContext1_stateSize;
  reg        [7:0]    SBox5Stage_tempContext1_stateID;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_0;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_1;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_2;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_3;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_4;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_5;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_6;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_7;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_8;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_9;
  reg        [254:0]  SBox5Stage_tempContext1_stateElements_10;
  reg        [254:0]  SBox5Stage_tempContext1_stateElement;
  wire                SBox5Stage_mulInput2_valid;
  wire       [254:0]  SBox5Stage_mulInput2_payload_op1;
  wire       [254:0]  SBox5Stage_mulInput2_payload_op2;
  wire                SBox5Stage_mul2Context_isFull;
  wire       [2:0]    SBox5Stage_mul2Context_fullRound;
  wire       [5:0]    SBox5Stage_mul2Context_partialRound;
  wire       [3:0]    SBox5Stage_mul2Context_stateIndex;
  wire       [3:0]    SBox5Stage_mul2Context_stateSize;
  wire       [7:0]    SBox5Stage_mul2Context_stateID;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_0;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_1;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_2;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_3;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_4;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_5;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_6;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_7;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_8;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_9;
  wire       [254:0]  SBox5Stage_mul2Context_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_1_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_1_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_1_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_1_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_1_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_1_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_1_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_2_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_2_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_2_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_2_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_2_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_2_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_2_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_3_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_3_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_3_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_3_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_3_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_3_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_3_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_4_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_4_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_4_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_4_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_4_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_4_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_4_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_5_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_5_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_5_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_5_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_5_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_5_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_5_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_6_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_6_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_6_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_6_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_6_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_6_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_6_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_7_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_7_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_7_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_7_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_7_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_7_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_7_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_8_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_8_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_8_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_8_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_8_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_8_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_8_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_9_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_9_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_9_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_9_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_9_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_9_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_9_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_10_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_10_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_10_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_10_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_10_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_10_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_10_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_11_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_11_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_11_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_11_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_11_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_11_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_11_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_12_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_12_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_12_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_12_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_12_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_12_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_12_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_13_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_13_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_13_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_13_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_13_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_13_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_13_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_14_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_14_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_14_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_14_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_14_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_14_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_14_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_15_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_15_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_15_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_15_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_15_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_15_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_15_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_16_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_16_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_16_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_16_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_16_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_16_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_16_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_17_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_17_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_17_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_17_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_17_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_17_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_17_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_18_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_18_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_18_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_18_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_18_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_18_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_18_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_19_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_19_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_19_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_19_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_19_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_19_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_19_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_20_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_20_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_20_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_20_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_20_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_20_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_20_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_21_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_21_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_21_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_21_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_21_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_21_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_21_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_22_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_22_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_22_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_22_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_22_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_22_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_22_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_23_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_23_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_23_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_23_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_23_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_23_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_23_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_24_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_24_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_24_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_24_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_24_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_24_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_24_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_25_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_25_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_25_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_25_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_25_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_25_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_25_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_26_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_26_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_26_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_26_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_26_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_26_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_26_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_27_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_27_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_27_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_27_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_27_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_27_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_27_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_28_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_28_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_28_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_28_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_28_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_28_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_28_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_29_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_29_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_29_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_29_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_29_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_29_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_29_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_30_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_30_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_30_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_30_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_30_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_30_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_30_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_31_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_31_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_31_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_31_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_31_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_31_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_31_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_32_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_32_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_32_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_32_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_32_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_32_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_32_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_33_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_33_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_33_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_33_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_33_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_33_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_33_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_34_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_34_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_34_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_34_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_34_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_34_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_34_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_35_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_35_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_35_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_35_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_35_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_35_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_35_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_36_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_36_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_36_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_36_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_36_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_36_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_36_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_37_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_37_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_37_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_37_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_37_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_37_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_37_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_38_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_38_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_38_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_38_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_38_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_38_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_38_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_39_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_39_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_39_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_39_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_39_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_39_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_39_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_40_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_40_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_40_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_40_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_40_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_40_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_40_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_41_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_41_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_41_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_41_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_41_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_41_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_41_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_42_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_42_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_42_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_42_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_42_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_42_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_42_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_43_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_43_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_43_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_43_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_43_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_43_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_43_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_44_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_44_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_44_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_44_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_44_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_44_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_44_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_45_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_45_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_45_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_45_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_45_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_45_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_45_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_46_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_46_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_46_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_46_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_46_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_46_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_46_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_47_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_47_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_47_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_47_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_47_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_47_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_47_stateElements_10;
  reg                 SBox5Stage_mul2Context_delay_48_isFull;
  reg        [2:0]    SBox5Stage_mul2Context_delay_48_fullRound;
  reg        [5:0]    SBox5Stage_mul2Context_delay_48_partialRound;
  reg        [3:0]    SBox5Stage_mul2Context_delay_48_stateIndex;
  reg        [3:0]    SBox5Stage_mul2Context_delay_48_stateSize;
  reg        [7:0]    SBox5Stage_mul2Context_delay_48_stateID;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_0;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_1;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_2;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_3;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_4;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_5;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_6;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_7;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_8;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_9;
  reg        [254:0]  SBox5Stage_mul2Context_delay_48_stateElements_10;
  reg                 SBox5Stage_tempContext2_isFull;
  reg        [2:0]    SBox5Stage_tempContext2_fullRound;
  reg        [5:0]    SBox5Stage_tempContext2_partialRound;
  reg        [3:0]    SBox5Stage_tempContext2_stateIndex;
  reg        [3:0]    SBox5Stage_tempContext2_stateSize;
  reg        [7:0]    SBox5Stage_tempContext2_stateID;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_0;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_1;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_2;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_3;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_4;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_5;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_6;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_7;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_8;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_9;
  reg        [254:0]  SBox5Stage_tempContext2_stateElements_10;
  wire                SBox5Stage_output_valid;
  wire                SBox5Stage_output_payload_isFull;
  wire       [2:0]    SBox5Stage_output_payload_fullRound;
  wire       [5:0]    SBox5Stage_output_payload_partialRound;
  wire       [3:0]    SBox5Stage_output_payload_stateIndex;
  wire       [3:0]    SBox5Stage_output_payload_stateSize;
  wire       [7:0]    SBox5Stage_output_payload_stateID;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_0;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_1;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_2;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_3;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_4;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_5;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_6;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_7;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_8;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_9;
  wire       [254:0]  SBox5Stage_output_payload_stateElements_10;
  wire       [254:0]  SBox5Stage_output_payload_stateElement;
  wire       [254:0]  AddRoundConstantStage_adderOperands_op1;
  wire       [254:0]  AddRoundConstantStage_adderOperands_op2;
  wire                AddRoundConstantStage_adderContext_isFull;
  wire       [2:0]    AddRoundConstantStage_adderContext_fullRound;
  wire       [5:0]    AddRoundConstantStage_adderContext_partialRound;
  wire       [3:0]    AddRoundConstantStage_adderContext_stateIndex;
  wire       [3:0]    AddRoundConstantStage_adderContext_stateSize;
  wire       [7:0]    AddRoundConstantStage_adderContext_stateID;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_0;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_1;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_2;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_3;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_4;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_5;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_6;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_7;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_8;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_9;
  wire       [254:0]  AddRoundConstantStage_adderContext_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_1_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_1_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_1_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_1_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_1_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_1_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_1_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_2_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_2_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_2_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_2_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_2_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_2_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_2_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_3_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_3_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_3_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_3_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_3_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_3_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_3_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_4_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_4_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_4_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_4_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_4_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_4_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_4_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_5_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_5_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_5_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_5_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_5_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_5_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_5_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_6_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_6_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_6_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_6_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_6_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_6_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_6_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_7_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_7_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_7_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_7_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_7_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_7_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_7_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_8_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_8_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_8_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_8_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_8_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_8_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_8_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_9_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_9_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_9_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_9_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_9_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_9_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_9_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_10_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_10_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_10_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_10_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_10_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_10_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_10_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_11_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_11_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_11_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_11_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_11_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_11_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_11_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_12_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_12_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_12_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_12_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_12_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_12_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_12_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_13_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_13_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_13_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_13_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_13_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_13_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_13_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_14_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_14_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_14_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_14_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_14_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_14_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_14_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_15_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_15_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_15_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_15_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_15_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_15_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_15_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_16_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_16_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_16_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_16_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_16_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_16_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_16_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_17_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_17_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_17_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_17_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_17_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_17_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_17_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_18_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_18_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_18_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_18_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_18_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_18_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_18_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_19_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_19_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_19_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_19_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_19_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_19_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_19_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_20_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_20_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_20_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_20_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_20_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_20_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_20_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_21_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_21_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_21_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_21_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_21_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_21_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_21_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_22_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_22_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_22_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_22_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_22_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_22_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_22_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_23_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_23_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_23_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_23_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_23_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_23_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_23_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_24_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_24_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_24_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_24_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_24_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_24_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_24_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_25_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_25_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_25_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_25_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_25_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_25_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_25_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_26_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_26_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_26_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_26_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_26_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_26_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_26_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_27_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_27_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_27_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_27_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_27_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_27_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_27_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_28_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_28_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_28_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_28_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_28_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_28_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_28_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_29_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_29_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_29_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_29_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_29_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_29_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_29_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_30_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_30_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_30_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_30_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_30_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_30_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_30_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_31_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_31_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_31_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_31_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_31_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_31_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_31_stateElements_10;
  reg                 AddRoundConstantStage_adderContext_delay_32_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContext_delay_32_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContext_delay_32_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_32_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContext_delay_32_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContext_delay_32_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContext_delay_32_stateElements_10;
  reg                 AddRoundConstantStage_adderContextDelayed_isFull;
  reg        [2:0]    AddRoundConstantStage_adderContextDelayed_fullRound;
  reg        [5:0]    AddRoundConstantStage_adderContextDelayed_partialRound;
  reg        [3:0]    AddRoundConstantStage_adderContextDelayed_stateIndex;
  reg        [3:0]    AddRoundConstantStage_adderContextDelayed_stateSize;
  reg        [7:0]    AddRoundConstantStage_adderContextDelayed_stateID;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_adderContextDelayed_stateElements_10;
  wire                AddRoundConstantStage_output_valid;
  wire                AddRoundConstantStage_output_payload_isFull;
  wire       [2:0]    AddRoundConstantStage_output_payload_fullRound;
  wire       [5:0]    AddRoundConstantStage_output_payload_partialRound;
  wire       [3:0]    AddRoundConstantStage_output_payload_stateIndex;
  wire       [3:0]    AddRoundConstantStage_output_payload_stateSize;
  wire       [7:0]    AddRoundConstantStage_output_payload_stateID;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_0;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_1;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_2;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_3;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_4;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_5;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_6;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_7;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_8;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_9;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElements_10;
  wire       [254:0]  AddRoundConstantStage_output_payload_stateElement;
  reg                 AddRoundConstantStage_output_regNext_valid;
  reg                 AddRoundConstantStage_output_regNext_payload_isFull;
  reg        [2:0]    AddRoundConstantStage_output_regNext_payload_fullRound;
  reg        [5:0]    AddRoundConstantStage_output_regNext_payload_partialRound;
  reg        [3:0]    AddRoundConstantStage_output_regNext_payload_stateIndex;
  reg        [3:0]    AddRoundConstantStage_output_regNext_payload_stateSize;
  reg        [7:0]    AddRoundConstantStage_output_regNext_payload_stateID;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_0;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_1;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_2;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_3;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_4;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_5;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_6;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_7;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_8;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_9;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElements_10;
  reg        [254:0]  AddRoundConstantStage_output_regNext_payload_stateElement;

  MontgomeryMultFlow SBox5Stage_montMultiplier0 (
    .io_input_valid           (SBox5Stage_mulInput0_valid                               ), //i
    .io_input_payload_op1     (SBox5Stage_mulInput0_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (SBox5Stage_mulInput0_payload_op2[254:0]                  ), //i
    .io_output_valid          (SBox5Stage_montMultiplier0_io_output_valid               ), //o
    .io_output_payload_res    (SBox5Stage_montMultiplier0_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                      ), //i
    .resetn                   (resetn                                                   )  //i
  );
  MontgomeryMultFlow SBox5Stage_montMultiplier1 (
    .io_input_valid           (SBox5Stage_mulInput1_valid                               ), //i
    .io_input_payload_op1     (SBox5Stage_mulInput1_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (SBox5Stage_mulInput1_payload_op2[254:0]                  ), //i
    .io_output_valid          (SBox5Stage_montMultiplier1_io_output_valid               ), //o
    .io_output_payload_res    (SBox5Stage_montMultiplier1_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                      ), //i
    .resetn                   (resetn                                                   )  //i
  );
  MontgomeryMultFlow SBox5Stage_montMultiplier2 (
    .io_input_valid           (SBox5Stage_mulInput2_valid                               ), //i
    .io_input_payload_op1     (SBox5Stage_mulInput2_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (SBox5Stage_mulInput2_payload_op2[254:0]                  ), //i
    .io_output_valid          (SBox5Stage_montMultiplier2_io_output_valid               ), //o
    .io_output_payload_res    (SBox5Stage_montMultiplier2_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                      ), //i
    .resetn                   (resetn                                                   )  //i
  );
  RoundConstantMem AddRoundConstantStage_constantMemory (
    .io_addr_isFull          (SBox5Stage_output_payload_isFull                     ), //i
    .io_addr_fullRound       (SBox5Stage_output_payload_fullRound[2:0]             ), //i
    .io_addr_partialRound    (SBox5Stage_output_payload_partialRound[5:0]          ), //i
    .io_addr_stateIndex      (SBox5Stage_output_payload_stateIndex[3:0]            ), //i
    .io_addr_stateSize       (SBox5Stage_output_payload_stateSize[3:0]             ), //i
    .io_data                 (AddRoundConstantStage_constantMemory_io_data[254:0]  )  //o
  );
  ModularAdderFlow AddRoundConstantStage_modAdder (
    .io_input_valid           (SBox5Stage_output_valid                                      ), //i
    .io_input_payload_op1     (AddRoundConstantStage_adderOperands_op1[254:0]               ), //i
    .io_input_payload_op2     (AddRoundConstantStage_adderOperands_op2[254:0]               ), //i
    .io_output_valid          (AddRoundConstantStage_modAdder_io_output_valid               ), //o
    .io_output_payload_res    (AddRoundConstantStage_modAdder_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                          ), //i
    .resetn                   (resetn                                                       )  //i
  );
  MDSMatrixMultiplier mDSMatrixMultiplier_1 (
    .io_input_valid                        (AddRoundConstantStage_output_regNext_valid                            ), //i
    .io_input_payload_isFull               (AddRoundConstantStage_output_regNext_payload_isFull                   ), //i
    .io_input_payload_fullRound            (AddRoundConstantStage_output_regNext_payload_fullRound[2:0]           ), //i
    .io_input_payload_partialRound         (AddRoundConstantStage_output_regNext_payload_partialRound[5:0]        ), //i
    .io_input_payload_stateIndex           (AddRoundConstantStage_output_regNext_payload_stateIndex[3:0]          ), //i
    .io_input_payload_stateSize            (AddRoundConstantStage_output_regNext_payload_stateSize[3:0]           ), //i
    .io_input_payload_stateID              (AddRoundConstantStage_output_regNext_payload_stateID[7:0]             ), //i
    .io_input_payload_stateElements_0      (AddRoundConstantStage_output_regNext_payload_stateElements_0[254:0]   ), //i
    .io_input_payload_stateElements_1      (AddRoundConstantStage_output_regNext_payload_stateElements_1[254:0]   ), //i
    .io_input_payload_stateElements_2      (AddRoundConstantStage_output_regNext_payload_stateElements_2[254:0]   ), //i
    .io_input_payload_stateElements_3      (AddRoundConstantStage_output_regNext_payload_stateElements_3[254:0]   ), //i
    .io_input_payload_stateElements_4      (AddRoundConstantStage_output_regNext_payload_stateElements_4[254:0]   ), //i
    .io_input_payload_stateElements_5      (AddRoundConstantStage_output_regNext_payload_stateElements_5[254:0]   ), //i
    .io_input_payload_stateElements_6      (AddRoundConstantStage_output_regNext_payload_stateElements_6[254:0]   ), //i
    .io_input_payload_stateElements_7      (AddRoundConstantStage_output_regNext_payload_stateElements_7[254:0]   ), //i
    .io_input_payload_stateElements_8      (AddRoundConstantStage_output_regNext_payload_stateElements_8[254:0]   ), //i
    .io_input_payload_stateElements_9      (AddRoundConstantStage_output_regNext_payload_stateElements_9[254:0]   ), //i
    .io_input_payload_stateElements_10     (AddRoundConstantStage_output_regNext_payload_stateElements_10[254:0]  ), //i
    .io_input_payload_stateElement         (AddRoundConstantStage_output_regNext_payload_stateElement[254:0]      ), //i
    .io_output_valid                       (mDSMatrixMultiplier_1_io_output_valid                                 ), //o
    .io_output_payload_isFull              (mDSMatrixMultiplier_1_io_output_payload_isFull                        ), //o
    .io_output_payload_fullRound           (mDSMatrixMultiplier_1_io_output_payload_fullRound[2:0]                ), //o
    .io_output_payload_partialRound        (mDSMatrixMultiplier_1_io_output_payload_partialRound[5:0]             ), //o
    .io_output_payload_stateSize           (mDSMatrixMultiplier_1_io_output_payload_stateSize[3:0]                ), //o
    .io_output_payload_stateID             (mDSMatrixMultiplier_1_io_output_payload_stateID[7:0]                  ), //o
    .io_output_payload_stateElements_0     (mDSMatrixMultiplier_1_io_output_payload_stateElements_0[254:0]        ), //o
    .io_output_payload_stateElements_1     (mDSMatrixMultiplier_1_io_output_payload_stateElements_1[254:0]        ), //o
    .io_output_payload_stateElements_2     (mDSMatrixMultiplier_1_io_output_payload_stateElements_2[254:0]        ), //o
    .io_output_payload_stateElements_3     (mDSMatrixMultiplier_1_io_output_payload_stateElements_3[254:0]        ), //o
    .io_output_payload_stateElements_4     (mDSMatrixMultiplier_1_io_output_payload_stateElements_4[254:0]        ), //o
    .io_output_payload_stateElements_5     (mDSMatrixMultiplier_1_io_output_payload_stateElements_5[254:0]        ), //o
    .io_output_payload_stateElements_6     (mDSMatrixMultiplier_1_io_output_payload_stateElements_6[254:0]        ), //o
    .io_output_payload_stateElements_7     (mDSMatrixMultiplier_1_io_output_payload_stateElements_7[254:0]        ), //o
    .io_output_payload_stateElements_8     (mDSMatrixMultiplier_1_io_output_payload_stateElements_8[254:0]        ), //o
    .io_output_payload_stateElements_9     (mDSMatrixMultiplier_1_io_output_payload_stateElements_9[254:0]        ), //o
    .io_output_payload_stateElements_10    (mDSMatrixMultiplier_1_io_output_payload_stateElements_10[254:0]       ), //o
    .io_output_payload_stateElements_11    (mDSMatrixMultiplier_1_io_output_payload_stateElements_11[254:0]       ), //o
    .clk                                   (clk                                                                   ), //i
    .resetn                                (resetn                                                                )  //i
  );
  MDSMatrixAdders mDSMatrixAdders_1 (
    .io_input_valid                        (mDSMatrixMultiplier_1_io_output_valid                            ), //i
    .io_input_payload_isFull               (mDSMatrixMultiplier_1_io_output_payload_isFull                   ), //i
    .io_input_payload_fullRound            (mDSMatrixMultiplier_1_io_output_payload_fullRound[2:0]           ), //i
    .io_input_payload_partialRound         (mDSMatrixMultiplier_1_io_output_payload_partialRound[5:0]        ), //i
    .io_input_payload_stateSize            (mDSMatrixMultiplier_1_io_output_payload_stateSize[3:0]           ), //i
    .io_input_payload_stateID              (mDSMatrixMultiplier_1_io_output_payload_stateID[7:0]             ), //i
    .io_input_payload_stateElements_0      (mDSMatrixMultiplier_1_io_output_payload_stateElements_0[254:0]   ), //i
    .io_input_payload_stateElements_1      (mDSMatrixMultiplier_1_io_output_payload_stateElements_1[254:0]   ), //i
    .io_input_payload_stateElements_2      (mDSMatrixMultiplier_1_io_output_payload_stateElements_2[254:0]   ), //i
    .io_input_payload_stateElements_3      (mDSMatrixMultiplier_1_io_output_payload_stateElements_3[254:0]   ), //i
    .io_input_payload_stateElements_4      (mDSMatrixMultiplier_1_io_output_payload_stateElements_4[254:0]   ), //i
    .io_input_payload_stateElements_5      (mDSMatrixMultiplier_1_io_output_payload_stateElements_5[254:0]   ), //i
    .io_input_payload_stateElements_6      (mDSMatrixMultiplier_1_io_output_payload_stateElements_6[254:0]   ), //i
    .io_input_payload_stateElements_7      (mDSMatrixMultiplier_1_io_output_payload_stateElements_7[254:0]   ), //i
    .io_input_payload_stateElements_8      (mDSMatrixMultiplier_1_io_output_payload_stateElements_8[254:0]   ), //i
    .io_input_payload_stateElements_9      (mDSMatrixMultiplier_1_io_output_payload_stateElements_9[254:0]   ), //i
    .io_input_payload_stateElements_10     (mDSMatrixMultiplier_1_io_output_payload_stateElements_10[254:0]  ), //i
    .io_input_payload_stateElements_11     (mDSMatrixMultiplier_1_io_output_payload_stateElements_11[254:0]  ), //i
    .io_output_valid                       (mDSMatrixAdders_1_io_output_valid                                ), //o
    .io_output_payload_isFull              (mDSMatrixAdders_1_io_output_payload_isFull                       ), //o
    .io_output_payload_fullRound           (mDSMatrixAdders_1_io_output_payload_fullRound[2:0]               ), //o
    .io_output_payload_partialRound        (mDSMatrixAdders_1_io_output_payload_partialRound[5:0]            ), //o
    .io_output_payload_stateSize           (mDSMatrixAdders_1_io_output_payload_stateSize[3:0]               ), //o
    .io_output_payload_stateID             (mDSMatrixAdders_1_io_output_payload_stateID[7:0]                 ), //o
    .io_output_payload_stateElements_0     (mDSMatrixAdders_1_io_output_payload_stateElements_0[254:0]       ), //o
    .io_output_payload_stateElements_1     (mDSMatrixAdders_1_io_output_payload_stateElements_1[254:0]       ), //o
    .io_output_payload_stateElements_2     (mDSMatrixAdders_1_io_output_payload_stateElements_2[254:0]       ), //o
    .io_output_payload_stateElements_3     (mDSMatrixAdders_1_io_output_payload_stateElements_3[254:0]       ), //o
    .io_output_payload_stateElements_4     (mDSMatrixAdders_1_io_output_payload_stateElements_4[254:0]       ), //o
    .io_output_payload_stateElements_5     (mDSMatrixAdders_1_io_output_payload_stateElements_5[254:0]       ), //o
    .io_output_payload_stateElements_6     (mDSMatrixAdders_1_io_output_payload_stateElements_6[254:0]       ), //o
    .io_output_payload_stateElements_7     (mDSMatrixAdders_1_io_output_payload_stateElements_7[254:0]       ), //o
    .io_output_payload_stateElements_8     (mDSMatrixAdders_1_io_output_payload_stateElements_8[254:0]       ), //o
    .io_output_payload_stateElements_9     (mDSMatrixAdders_1_io_output_payload_stateElements_9[254:0]       ), //o
    .io_output_payload_stateElements_10    (mDSMatrixAdders_1_io_output_payload_stateElements_10[254:0]      ), //o
    .io_output_payload_stateElements_11    (mDSMatrixAdders_1_io_output_payload_stateElements_11[254:0]      ), //o
    .clk                                   (clk                                                              ), //i
    .resetn                                (resetn                                                           )  //i
  );
  assign SBox5Stage_mulInput0_valid = io_input_valid;
  assign SBox5Stage_mulInput0_payload_op1 = io_input_payload_stateElement;
  assign SBox5Stage_mulInput0_payload_op2 = io_input_payload_stateElement;
  assign SBox5Stage_mulInput1_valid = SBox5Stage_montMultiplier0_io_output_valid;
  assign SBox5Stage_mulInput1_payload_op1 = SBox5Stage_montMultiplier0_io_output_payload_res;
  assign SBox5Stage_mulInput1_payload_op2 = SBox5Stage_montMultiplier0_io_output_payload_res;
  assign SBox5Stage_mulInput2_valid = SBox5Stage_montMultiplier1_io_output_valid;
  assign SBox5Stage_mulInput2_payload_op1 = SBox5Stage_montMultiplier1_io_output_payload_res;
  assign SBox5Stage_mulInput2_payload_op2 = SBox5Stage_tempContext1_stateElement;
  assign SBox5Stage_mul2Context_isFull = SBox5Stage_tempContext1_isFull;
  assign SBox5Stage_mul2Context_fullRound = SBox5Stage_tempContext1_fullRound;
  assign SBox5Stage_mul2Context_partialRound = SBox5Stage_tempContext1_partialRound;
  assign SBox5Stage_mul2Context_stateIndex = SBox5Stage_tempContext1_stateIndex;
  assign SBox5Stage_mul2Context_stateSize = SBox5Stage_tempContext1_stateSize;
  assign SBox5Stage_mul2Context_stateID = SBox5Stage_tempContext1_stateID;
  assign SBox5Stage_mul2Context_stateElements_0 = SBox5Stage_tempContext1_stateElements_0;
  assign SBox5Stage_mul2Context_stateElements_1 = SBox5Stage_tempContext1_stateElements_1;
  assign SBox5Stage_mul2Context_stateElements_2 = SBox5Stage_tempContext1_stateElements_2;
  assign SBox5Stage_mul2Context_stateElements_3 = SBox5Stage_tempContext1_stateElements_3;
  assign SBox5Stage_mul2Context_stateElements_4 = SBox5Stage_tempContext1_stateElements_4;
  assign SBox5Stage_mul2Context_stateElements_5 = SBox5Stage_tempContext1_stateElements_5;
  assign SBox5Stage_mul2Context_stateElements_6 = SBox5Stage_tempContext1_stateElements_6;
  assign SBox5Stage_mul2Context_stateElements_7 = SBox5Stage_tempContext1_stateElements_7;
  assign SBox5Stage_mul2Context_stateElements_8 = SBox5Stage_tempContext1_stateElements_8;
  assign SBox5Stage_mul2Context_stateElements_9 = SBox5Stage_tempContext1_stateElements_9;
  assign SBox5Stage_mul2Context_stateElements_10 = SBox5Stage_tempContext1_stateElements_10;
  assign SBox5Stage_output_valid = SBox5Stage_montMultiplier2_io_output_valid;
  assign SBox5Stage_output_payload_isFull = SBox5Stage_tempContext2_isFull;
  assign SBox5Stage_output_payload_fullRound = SBox5Stage_tempContext2_fullRound;
  assign SBox5Stage_output_payload_partialRound = SBox5Stage_tempContext2_partialRound;
  assign SBox5Stage_output_payload_stateIndex = SBox5Stage_tempContext2_stateIndex;
  assign SBox5Stage_output_payload_stateSize = SBox5Stage_tempContext2_stateSize;
  assign SBox5Stage_output_payload_stateID = SBox5Stage_tempContext2_stateID;
  assign SBox5Stage_output_payload_stateElements_0 = SBox5Stage_tempContext2_stateElements_0;
  assign SBox5Stage_output_payload_stateElements_1 = SBox5Stage_tempContext2_stateElements_1;
  assign SBox5Stage_output_payload_stateElements_2 = SBox5Stage_tempContext2_stateElements_2;
  assign SBox5Stage_output_payload_stateElements_3 = SBox5Stage_tempContext2_stateElements_3;
  assign SBox5Stage_output_payload_stateElements_4 = SBox5Stage_tempContext2_stateElements_4;
  assign SBox5Stage_output_payload_stateElements_5 = SBox5Stage_tempContext2_stateElements_5;
  assign SBox5Stage_output_payload_stateElements_6 = SBox5Stage_tempContext2_stateElements_6;
  assign SBox5Stage_output_payload_stateElements_7 = SBox5Stage_tempContext2_stateElements_7;
  assign SBox5Stage_output_payload_stateElements_8 = SBox5Stage_tempContext2_stateElements_8;
  assign SBox5Stage_output_payload_stateElements_9 = SBox5Stage_tempContext2_stateElements_9;
  assign SBox5Stage_output_payload_stateElements_10 = SBox5Stage_tempContext2_stateElements_10;
  assign SBox5Stage_output_payload_stateElement = SBox5Stage_montMultiplier2_io_output_payload_res;
  assign AddRoundConstantStage_adderOperands_op1 = SBox5Stage_output_payload_stateElement;
  assign AddRoundConstantStage_adderOperands_op2 = AddRoundConstantStage_constantMemory_io_data;
  assign AddRoundConstantStage_adderContext_isFull = SBox5Stage_output_payload_isFull;
  assign AddRoundConstantStage_adderContext_fullRound = SBox5Stage_output_payload_fullRound;
  assign AddRoundConstantStage_adderContext_partialRound = SBox5Stage_output_payload_partialRound;
  assign AddRoundConstantStage_adderContext_stateIndex = SBox5Stage_output_payload_stateIndex;
  assign AddRoundConstantStage_adderContext_stateSize = SBox5Stage_output_payload_stateSize;
  assign AddRoundConstantStage_adderContext_stateID = SBox5Stage_output_payload_stateID;
  assign AddRoundConstantStage_adderContext_stateElements_0 = SBox5Stage_output_payload_stateElements_0;
  assign AddRoundConstantStage_adderContext_stateElements_1 = SBox5Stage_output_payload_stateElements_1;
  assign AddRoundConstantStage_adderContext_stateElements_2 = SBox5Stage_output_payload_stateElements_2;
  assign AddRoundConstantStage_adderContext_stateElements_3 = SBox5Stage_output_payload_stateElements_3;
  assign AddRoundConstantStage_adderContext_stateElements_4 = SBox5Stage_output_payload_stateElements_4;
  assign AddRoundConstantStage_adderContext_stateElements_5 = SBox5Stage_output_payload_stateElements_5;
  assign AddRoundConstantStage_adderContext_stateElements_6 = SBox5Stage_output_payload_stateElements_6;
  assign AddRoundConstantStage_adderContext_stateElements_7 = SBox5Stage_output_payload_stateElements_7;
  assign AddRoundConstantStage_adderContext_stateElements_8 = SBox5Stage_output_payload_stateElements_8;
  assign AddRoundConstantStage_adderContext_stateElements_9 = SBox5Stage_output_payload_stateElements_9;
  assign AddRoundConstantStage_adderContext_stateElements_10 = SBox5Stage_output_payload_stateElements_10;
  assign AddRoundConstantStage_output_valid = AddRoundConstantStage_modAdder_io_output_valid;
  assign AddRoundConstantStage_output_payload_isFull = AddRoundConstantStage_adderContextDelayed_isFull;
  assign AddRoundConstantStage_output_payload_fullRound = AddRoundConstantStage_adderContextDelayed_fullRound;
  assign AddRoundConstantStage_output_payload_partialRound = AddRoundConstantStage_adderContextDelayed_partialRound;
  assign AddRoundConstantStage_output_payload_stateIndex = AddRoundConstantStage_adderContextDelayed_stateIndex;
  assign AddRoundConstantStage_output_payload_stateSize = AddRoundConstantStage_adderContextDelayed_stateSize;
  assign AddRoundConstantStage_output_payload_stateID = AddRoundConstantStage_adderContextDelayed_stateID;
  assign AddRoundConstantStage_output_payload_stateElements_0 = AddRoundConstantStage_adderContextDelayed_stateElements_0;
  assign AddRoundConstantStage_output_payload_stateElements_1 = AddRoundConstantStage_adderContextDelayed_stateElements_1;
  assign AddRoundConstantStage_output_payload_stateElements_2 = AddRoundConstantStage_adderContextDelayed_stateElements_2;
  assign AddRoundConstantStage_output_payload_stateElements_3 = AddRoundConstantStage_adderContextDelayed_stateElements_3;
  assign AddRoundConstantStage_output_payload_stateElements_4 = AddRoundConstantStage_adderContextDelayed_stateElements_4;
  assign AddRoundConstantStage_output_payload_stateElements_5 = AddRoundConstantStage_adderContextDelayed_stateElements_5;
  assign AddRoundConstantStage_output_payload_stateElements_6 = AddRoundConstantStage_adderContextDelayed_stateElements_6;
  assign AddRoundConstantStage_output_payload_stateElements_7 = AddRoundConstantStage_adderContextDelayed_stateElements_7;
  assign AddRoundConstantStage_output_payload_stateElements_8 = AddRoundConstantStage_adderContextDelayed_stateElements_8;
  assign AddRoundConstantStage_output_payload_stateElements_9 = AddRoundConstantStage_adderContextDelayed_stateElements_9;
  assign AddRoundConstantStage_output_payload_stateElements_10 = AddRoundConstantStage_adderContextDelayed_stateElements_10;
  assign AddRoundConstantStage_output_payload_stateElement = AddRoundConstantStage_modAdder_io_output_payload_res;
  assign io_output_valid = mDSMatrixAdders_1_io_output_valid;
  assign io_output_payload_isFull = mDSMatrixAdders_1_io_output_payload_isFull;
  assign io_output_payload_fullRound = mDSMatrixAdders_1_io_output_payload_fullRound;
  assign io_output_payload_partialRound = mDSMatrixAdders_1_io_output_payload_partialRound;
  assign io_output_payload_stateSize = mDSMatrixAdders_1_io_output_payload_stateSize;
  assign io_output_payload_stateID = mDSMatrixAdders_1_io_output_payload_stateID;
  assign io_output_payload_stateElements_0 = mDSMatrixAdders_1_io_output_payload_stateElements_0;
  assign io_output_payload_stateElements_1 = mDSMatrixAdders_1_io_output_payload_stateElements_1;
  assign io_output_payload_stateElements_2 = mDSMatrixAdders_1_io_output_payload_stateElements_2;
  assign io_output_payload_stateElements_3 = mDSMatrixAdders_1_io_output_payload_stateElements_3;
  assign io_output_payload_stateElements_4 = mDSMatrixAdders_1_io_output_payload_stateElements_4;
  assign io_output_payload_stateElements_5 = mDSMatrixAdders_1_io_output_payload_stateElements_5;
  assign io_output_payload_stateElements_6 = mDSMatrixAdders_1_io_output_payload_stateElements_6;
  assign io_output_payload_stateElements_7 = mDSMatrixAdders_1_io_output_payload_stateElements_7;
  assign io_output_payload_stateElements_8 = mDSMatrixAdders_1_io_output_payload_stateElements_8;
  assign io_output_payload_stateElements_9 = mDSMatrixAdders_1_io_output_payload_stateElements_9;
  assign io_output_payload_stateElements_10 = mDSMatrixAdders_1_io_output_payload_stateElements_10;
  assign io_output_payload_stateElements_11 = mDSMatrixAdders_1_io_output_payload_stateElements_11;
  always @(posedge clk) begin
    io_input_payload_delay_1_isFull <= io_input_payload_isFull;
    io_input_payload_delay_1_fullRound <= io_input_payload_fullRound;
    io_input_payload_delay_1_partialRound <= io_input_payload_partialRound;
    io_input_payload_delay_1_stateIndex <= io_input_payload_stateIndex;
    io_input_payload_delay_1_stateSize <= io_input_payload_stateSize;
    io_input_payload_delay_1_stateID <= io_input_payload_stateID;
    io_input_payload_delay_1_stateElements_0 <= io_input_payload_stateElements_0;
    io_input_payload_delay_1_stateElements_1 <= io_input_payload_stateElements_1;
    io_input_payload_delay_1_stateElements_2 <= io_input_payload_stateElements_2;
    io_input_payload_delay_1_stateElements_3 <= io_input_payload_stateElements_3;
    io_input_payload_delay_1_stateElements_4 <= io_input_payload_stateElements_4;
    io_input_payload_delay_1_stateElements_5 <= io_input_payload_stateElements_5;
    io_input_payload_delay_1_stateElements_6 <= io_input_payload_stateElements_6;
    io_input_payload_delay_1_stateElements_7 <= io_input_payload_stateElements_7;
    io_input_payload_delay_1_stateElements_8 <= io_input_payload_stateElements_8;
    io_input_payload_delay_1_stateElements_9 <= io_input_payload_stateElements_9;
    io_input_payload_delay_1_stateElements_10 <= io_input_payload_stateElements_10;
    io_input_payload_delay_1_stateElement <= io_input_payload_stateElement;
    io_input_payload_delay_2_isFull <= io_input_payload_delay_1_isFull;
    io_input_payload_delay_2_fullRound <= io_input_payload_delay_1_fullRound;
    io_input_payload_delay_2_partialRound <= io_input_payload_delay_1_partialRound;
    io_input_payload_delay_2_stateIndex <= io_input_payload_delay_1_stateIndex;
    io_input_payload_delay_2_stateSize <= io_input_payload_delay_1_stateSize;
    io_input_payload_delay_2_stateID <= io_input_payload_delay_1_stateID;
    io_input_payload_delay_2_stateElements_0 <= io_input_payload_delay_1_stateElements_0;
    io_input_payload_delay_2_stateElements_1 <= io_input_payload_delay_1_stateElements_1;
    io_input_payload_delay_2_stateElements_2 <= io_input_payload_delay_1_stateElements_2;
    io_input_payload_delay_2_stateElements_3 <= io_input_payload_delay_1_stateElements_3;
    io_input_payload_delay_2_stateElements_4 <= io_input_payload_delay_1_stateElements_4;
    io_input_payload_delay_2_stateElements_5 <= io_input_payload_delay_1_stateElements_5;
    io_input_payload_delay_2_stateElements_6 <= io_input_payload_delay_1_stateElements_6;
    io_input_payload_delay_2_stateElements_7 <= io_input_payload_delay_1_stateElements_7;
    io_input_payload_delay_2_stateElements_8 <= io_input_payload_delay_1_stateElements_8;
    io_input_payload_delay_2_stateElements_9 <= io_input_payload_delay_1_stateElements_9;
    io_input_payload_delay_2_stateElements_10 <= io_input_payload_delay_1_stateElements_10;
    io_input_payload_delay_2_stateElement <= io_input_payload_delay_1_stateElement;
    io_input_payload_delay_3_isFull <= io_input_payload_delay_2_isFull;
    io_input_payload_delay_3_fullRound <= io_input_payload_delay_2_fullRound;
    io_input_payload_delay_3_partialRound <= io_input_payload_delay_2_partialRound;
    io_input_payload_delay_3_stateIndex <= io_input_payload_delay_2_stateIndex;
    io_input_payload_delay_3_stateSize <= io_input_payload_delay_2_stateSize;
    io_input_payload_delay_3_stateID <= io_input_payload_delay_2_stateID;
    io_input_payload_delay_3_stateElements_0 <= io_input_payload_delay_2_stateElements_0;
    io_input_payload_delay_3_stateElements_1 <= io_input_payload_delay_2_stateElements_1;
    io_input_payload_delay_3_stateElements_2 <= io_input_payload_delay_2_stateElements_2;
    io_input_payload_delay_3_stateElements_3 <= io_input_payload_delay_2_stateElements_3;
    io_input_payload_delay_3_stateElements_4 <= io_input_payload_delay_2_stateElements_4;
    io_input_payload_delay_3_stateElements_5 <= io_input_payload_delay_2_stateElements_5;
    io_input_payload_delay_3_stateElements_6 <= io_input_payload_delay_2_stateElements_6;
    io_input_payload_delay_3_stateElements_7 <= io_input_payload_delay_2_stateElements_7;
    io_input_payload_delay_3_stateElements_8 <= io_input_payload_delay_2_stateElements_8;
    io_input_payload_delay_3_stateElements_9 <= io_input_payload_delay_2_stateElements_9;
    io_input_payload_delay_3_stateElements_10 <= io_input_payload_delay_2_stateElements_10;
    io_input_payload_delay_3_stateElement <= io_input_payload_delay_2_stateElement;
    io_input_payload_delay_4_isFull <= io_input_payload_delay_3_isFull;
    io_input_payload_delay_4_fullRound <= io_input_payload_delay_3_fullRound;
    io_input_payload_delay_4_partialRound <= io_input_payload_delay_3_partialRound;
    io_input_payload_delay_4_stateIndex <= io_input_payload_delay_3_stateIndex;
    io_input_payload_delay_4_stateSize <= io_input_payload_delay_3_stateSize;
    io_input_payload_delay_4_stateID <= io_input_payload_delay_3_stateID;
    io_input_payload_delay_4_stateElements_0 <= io_input_payload_delay_3_stateElements_0;
    io_input_payload_delay_4_stateElements_1 <= io_input_payload_delay_3_stateElements_1;
    io_input_payload_delay_4_stateElements_2 <= io_input_payload_delay_3_stateElements_2;
    io_input_payload_delay_4_stateElements_3 <= io_input_payload_delay_3_stateElements_3;
    io_input_payload_delay_4_stateElements_4 <= io_input_payload_delay_3_stateElements_4;
    io_input_payload_delay_4_stateElements_5 <= io_input_payload_delay_3_stateElements_5;
    io_input_payload_delay_4_stateElements_6 <= io_input_payload_delay_3_stateElements_6;
    io_input_payload_delay_4_stateElements_7 <= io_input_payload_delay_3_stateElements_7;
    io_input_payload_delay_4_stateElements_8 <= io_input_payload_delay_3_stateElements_8;
    io_input_payload_delay_4_stateElements_9 <= io_input_payload_delay_3_stateElements_9;
    io_input_payload_delay_4_stateElements_10 <= io_input_payload_delay_3_stateElements_10;
    io_input_payload_delay_4_stateElement <= io_input_payload_delay_3_stateElement;
    io_input_payload_delay_5_isFull <= io_input_payload_delay_4_isFull;
    io_input_payload_delay_5_fullRound <= io_input_payload_delay_4_fullRound;
    io_input_payload_delay_5_partialRound <= io_input_payload_delay_4_partialRound;
    io_input_payload_delay_5_stateIndex <= io_input_payload_delay_4_stateIndex;
    io_input_payload_delay_5_stateSize <= io_input_payload_delay_4_stateSize;
    io_input_payload_delay_5_stateID <= io_input_payload_delay_4_stateID;
    io_input_payload_delay_5_stateElements_0 <= io_input_payload_delay_4_stateElements_0;
    io_input_payload_delay_5_stateElements_1 <= io_input_payload_delay_4_stateElements_1;
    io_input_payload_delay_5_stateElements_2 <= io_input_payload_delay_4_stateElements_2;
    io_input_payload_delay_5_stateElements_3 <= io_input_payload_delay_4_stateElements_3;
    io_input_payload_delay_5_stateElements_4 <= io_input_payload_delay_4_stateElements_4;
    io_input_payload_delay_5_stateElements_5 <= io_input_payload_delay_4_stateElements_5;
    io_input_payload_delay_5_stateElements_6 <= io_input_payload_delay_4_stateElements_6;
    io_input_payload_delay_5_stateElements_7 <= io_input_payload_delay_4_stateElements_7;
    io_input_payload_delay_5_stateElements_8 <= io_input_payload_delay_4_stateElements_8;
    io_input_payload_delay_5_stateElements_9 <= io_input_payload_delay_4_stateElements_9;
    io_input_payload_delay_5_stateElements_10 <= io_input_payload_delay_4_stateElements_10;
    io_input_payload_delay_5_stateElement <= io_input_payload_delay_4_stateElement;
    io_input_payload_delay_6_isFull <= io_input_payload_delay_5_isFull;
    io_input_payload_delay_6_fullRound <= io_input_payload_delay_5_fullRound;
    io_input_payload_delay_6_partialRound <= io_input_payload_delay_5_partialRound;
    io_input_payload_delay_6_stateIndex <= io_input_payload_delay_5_stateIndex;
    io_input_payload_delay_6_stateSize <= io_input_payload_delay_5_stateSize;
    io_input_payload_delay_6_stateID <= io_input_payload_delay_5_stateID;
    io_input_payload_delay_6_stateElements_0 <= io_input_payload_delay_5_stateElements_0;
    io_input_payload_delay_6_stateElements_1 <= io_input_payload_delay_5_stateElements_1;
    io_input_payload_delay_6_stateElements_2 <= io_input_payload_delay_5_stateElements_2;
    io_input_payload_delay_6_stateElements_3 <= io_input_payload_delay_5_stateElements_3;
    io_input_payload_delay_6_stateElements_4 <= io_input_payload_delay_5_stateElements_4;
    io_input_payload_delay_6_stateElements_5 <= io_input_payload_delay_5_stateElements_5;
    io_input_payload_delay_6_stateElements_6 <= io_input_payload_delay_5_stateElements_6;
    io_input_payload_delay_6_stateElements_7 <= io_input_payload_delay_5_stateElements_7;
    io_input_payload_delay_6_stateElements_8 <= io_input_payload_delay_5_stateElements_8;
    io_input_payload_delay_6_stateElements_9 <= io_input_payload_delay_5_stateElements_9;
    io_input_payload_delay_6_stateElements_10 <= io_input_payload_delay_5_stateElements_10;
    io_input_payload_delay_6_stateElement <= io_input_payload_delay_5_stateElement;
    io_input_payload_delay_7_isFull <= io_input_payload_delay_6_isFull;
    io_input_payload_delay_7_fullRound <= io_input_payload_delay_6_fullRound;
    io_input_payload_delay_7_partialRound <= io_input_payload_delay_6_partialRound;
    io_input_payload_delay_7_stateIndex <= io_input_payload_delay_6_stateIndex;
    io_input_payload_delay_7_stateSize <= io_input_payload_delay_6_stateSize;
    io_input_payload_delay_7_stateID <= io_input_payload_delay_6_stateID;
    io_input_payload_delay_7_stateElements_0 <= io_input_payload_delay_6_stateElements_0;
    io_input_payload_delay_7_stateElements_1 <= io_input_payload_delay_6_stateElements_1;
    io_input_payload_delay_7_stateElements_2 <= io_input_payload_delay_6_stateElements_2;
    io_input_payload_delay_7_stateElements_3 <= io_input_payload_delay_6_stateElements_3;
    io_input_payload_delay_7_stateElements_4 <= io_input_payload_delay_6_stateElements_4;
    io_input_payload_delay_7_stateElements_5 <= io_input_payload_delay_6_stateElements_5;
    io_input_payload_delay_7_stateElements_6 <= io_input_payload_delay_6_stateElements_6;
    io_input_payload_delay_7_stateElements_7 <= io_input_payload_delay_6_stateElements_7;
    io_input_payload_delay_7_stateElements_8 <= io_input_payload_delay_6_stateElements_8;
    io_input_payload_delay_7_stateElements_9 <= io_input_payload_delay_6_stateElements_9;
    io_input_payload_delay_7_stateElements_10 <= io_input_payload_delay_6_stateElements_10;
    io_input_payload_delay_7_stateElement <= io_input_payload_delay_6_stateElement;
    io_input_payload_delay_8_isFull <= io_input_payload_delay_7_isFull;
    io_input_payload_delay_8_fullRound <= io_input_payload_delay_7_fullRound;
    io_input_payload_delay_8_partialRound <= io_input_payload_delay_7_partialRound;
    io_input_payload_delay_8_stateIndex <= io_input_payload_delay_7_stateIndex;
    io_input_payload_delay_8_stateSize <= io_input_payload_delay_7_stateSize;
    io_input_payload_delay_8_stateID <= io_input_payload_delay_7_stateID;
    io_input_payload_delay_8_stateElements_0 <= io_input_payload_delay_7_stateElements_0;
    io_input_payload_delay_8_stateElements_1 <= io_input_payload_delay_7_stateElements_1;
    io_input_payload_delay_8_stateElements_2 <= io_input_payload_delay_7_stateElements_2;
    io_input_payload_delay_8_stateElements_3 <= io_input_payload_delay_7_stateElements_3;
    io_input_payload_delay_8_stateElements_4 <= io_input_payload_delay_7_stateElements_4;
    io_input_payload_delay_8_stateElements_5 <= io_input_payload_delay_7_stateElements_5;
    io_input_payload_delay_8_stateElements_6 <= io_input_payload_delay_7_stateElements_6;
    io_input_payload_delay_8_stateElements_7 <= io_input_payload_delay_7_stateElements_7;
    io_input_payload_delay_8_stateElements_8 <= io_input_payload_delay_7_stateElements_8;
    io_input_payload_delay_8_stateElements_9 <= io_input_payload_delay_7_stateElements_9;
    io_input_payload_delay_8_stateElements_10 <= io_input_payload_delay_7_stateElements_10;
    io_input_payload_delay_8_stateElement <= io_input_payload_delay_7_stateElement;
    io_input_payload_delay_9_isFull <= io_input_payload_delay_8_isFull;
    io_input_payload_delay_9_fullRound <= io_input_payload_delay_8_fullRound;
    io_input_payload_delay_9_partialRound <= io_input_payload_delay_8_partialRound;
    io_input_payload_delay_9_stateIndex <= io_input_payload_delay_8_stateIndex;
    io_input_payload_delay_9_stateSize <= io_input_payload_delay_8_stateSize;
    io_input_payload_delay_9_stateID <= io_input_payload_delay_8_stateID;
    io_input_payload_delay_9_stateElements_0 <= io_input_payload_delay_8_stateElements_0;
    io_input_payload_delay_9_stateElements_1 <= io_input_payload_delay_8_stateElements_1;
    io_input_payload_delay_9_stateElements_2 <= io_input_payload_delay_8_stateElements_2;
    io_input_payload_delay_9_stateElements_3 <= io_input_payload_delay_8_stateElements_3;
    io_input_payload_delay_9_stateElements_4 <= io_input_payload_delay_8_stateElements_4;
    io_input_payload_delay_9_stateElements_5 <= io_input_payload_delay_8_stateElements_5;
    io_input_payload_delay_9_stateElements_6 <= io_input_payload_delay_8_stateElements_6;
    io_input_payload_delay_9_stateElements_7 <= io_input_payload_delay_8_stateElements_7;
    io_input_payload_delay_9_stateElements_8 <= io_input_payload_delay_8_stateElements_8;
    io_input_payload_delay_9_stateElements_9 <= io_input_payload_delay_8_stateElements_9;
    io_input_payload_delay_9_stateElements_10 <= io_input_payload_delay_8_stateElements_10;
    io_input_payload_delay_9_stateElement <= io_input_payload_delay_8_stateElement;
    io_input_payload_delay_10_isFull <= io_input_payload_delay_9_isFull;
    io_input_payload_delay_10_fullRound <= io_input_payload_delay_9_fullRound;
    io_input_payload_delay_10_partialRound <= io_input_payload_delay_9_partialRound;
    io_input_payload_delay_10_stateIndex <= io_input_payload_delay_9_stateIndex;
    io_input_payload_delay_10_stateSize <= io_input_payload_delay_9_stateSize;
    io_input_payload_delay_10_stateID <= io_input_payload_delay_9_stateID;
    io_input_payload_delay_10_stateElements_0 <= io_input_payload_delay_9_stateElements_0;
    io_input_payload_delay_10_stateElements_1 <= io_input_payload_delay_9_stateElements_1;
    io_input_payload_delay_10_stateElements_2 <= io_input_payload_delay_9_stateElements_2;
    io_input_payload_delay_10_stateElements_3 <= io_input_payload_delay_9_stateElements_3;
    io_input_payload_delay_10_stateElements_4 <= io_input_payload_delay_9_stateElements_4;
    io_input_payload_delay_10_stateElements_5 <= io_input_payload_delay_9_stateElements_5;
    io_input_payload_delay_10_stateElements_6 <= io_input_payload_delay_9_stateElements_6;
    io_input_payload_delay_10_stateElements_7 <= io_input_payload_delay_9_stateElements_7;
    io_input_payload_delay_10_stateElements_8 <= io_input_payload_delay_9_stateElements_8;
    io_input_payload_delay_10_stateElements_9 <= io_input_payload_delay_9_stateElements_9;
    io_input_payload_delay_10_stateElements_10 <= io_input_payload_delay_9_stateElements_10;
    io_input_payload_delay_10_stateElement <= io_input_payload_delay_9_stateElement;
    io_input_payload_delay_11_isFull <= io_input_payload_delay_10_isFull;
    io_input_payload_delay_11_fullRound <= io_input_payload_delay_10_fullRound;
    io_input_payload_delay_11_partialRound <= io_input_payload_delay_10_partialRound;
    io_input_payload_delay_11_stateIndex <= io_input_payload_delay_10_stateIndex;
    io_input_payload_delay_11_stateSize <= io_input_payload_delay_10_stateSize;
    io_input_payload_delay_11_stateID <= io_input_payload_delay_10_stateID;
    io_input_payload_delay_11_stateElements_0 <= io_input_payload_delay_10_stateElements_0;
    io_input_payload_delay_11_stateElements_1 <= io_input_payload_delay_10_stateElements_1;
    io_input_payload_delay_11_stateElements_2 <= io_input_payload_delay_10_stateElements_2;
    io_input_payload_delay_11_stateElements_3 <= io_input_payload_delay_10_stateElements_3;
    io_input_payload_delay_11_stateElements_4 <= io_input_payload_delay_10_stateElements_4;
    io_input_payload_delay_11_stateElements_5 <= io_input_payload_delay_10_stateElements_5;
    io_input_payload_delay_11_stateElements_6 <= io_input_payload_delay_10_stateElements_6;
    io_input_payload_delay_11_stateElements_7 <= io_input_payload_delay_10_stateElements_7;
    io_input_payload_delay_11_stateElements_8 <= io_input_payload_delay_10_stateElements_8;
    io_input_payload_delay_11_stateElements_9 <= io_input_payload_delay_10_stateElements_9;
    io_input_payload_delay_11_stateElements_10 <= io_input_payload_delay_10_stateElements_10;
    io_input_payload_delay_11_stateElement <= io_input_payload_delay_10_stateElement;
    io_input_payload_delay_12_isFull <= io_input_payload_delay_11_isFull;
    io_input_payload_delay_12_fullRound <= io_input_payload_delay_11_fullRound;
    io_input_payload_delay_12_partialRound <= io_input_payload_delay_11_partialRound;
    io_input_payload_delay_12_stateIndex <= io_input_payload_delay_11_stateIndex;
    io_input_payload_delay_12_stateSize <= io_input_payload_delay_11_stateSize;
    io_input_payload_delay_12_stateID <= io_input_payload_delay_11_stateID;
    io_input_payload_delay_12_stateElements_0 <= io_input_payload_delay_11_stateElements_0;
    io_input_payload_delay_12_stateElements_1 <= io_input_payload_delay_11_stateElements_1;
    io_input_payload_delay_12_stateElements_2 <= io_input_payload_delay_11_stateElements_2;
    io_input_payload_delay_12_stateElements_3 <= io_input_payload_delay_11_stateElements_3;
    io_input_payload_delay_12_stateElements_4 <= io_input_payload_delay_11_stateElements_4;
    io_input_payload_delay_12_stateElements_5 <= io_input_payload_delay_11_stateElements_5;
    io_input_payload_delay_12_stateElements_6 <= io_input_payload_delay_11_stateElements_6;
    io_input_payload_delay_12_stateElements_7 <= io_input_payload_delay_11_stateElements_7;
    io_input_payload_delay_12_stateElements_8 <= io_input_payload_delay_11_stateElements_8;
    io_input_payload_delay_12_stateElements_9 <= io_input_payload_delay_11_stateElements_9;
    io_input_payload_delay_12_stateElements_10 <= io_input_payload_delay_11_stateElements_10;
    io_input_payload_delay_12_stateElement <= io_input_payload_delay_11_stateElement;
    io_input_payload_delay_13_isFull <= io_input_payload_delay_12_isFull;
    io_input_payload_delay_13_fullRound <= io_input_payload_delay_12_fullRound;
    io_input_payload_delay_13_partialRound <= io_input_payload_delay_12_partialRound;
    io_input_payload_delay_13_stateIndex <= io_input_payload_delay_12_stateIndex;
    io_input_payload_delay_13_stateSize <= io_input_payload_delay_12_stateSize;
    io_input_payload_delay_13_stateID <= io_input_payload_delay_12_stateID;
    io_input_payload_delay_13_stateElements_0 <= io_input_payload_delay_12_stateElements_0;
    io_input_payload_delay_13_stateElements_1 <= io_input_payload_delay_12_stateElements_1;
    io_input_payload_delay_13_stateElements_2 <= io_input_payload_delay_12_stateElements_2;
    io_input_payload_delay_13_stateElements_3 <= io_input_payload_delay_12_stateElements_3;
    io_input_payload_delay_13_stateElements_4 <= io_input_payload_delay_12_stateElements_4;
    io_input_payload_delay_13_stateElements_5 <= io_input_payload_delay_12_stateElements_5;
    io_input_payload_delay_13_stateElements_6 <= io_input_payload_delay_12_stateElements_6;
    io_input_payload_delay_13_stateElements_7 <= io_input_payload_delay_12_stateElements_7;
    io_input_payload_delay_13_stateElements_8 <= io_input_payload_delay_12_stateElements_8;
    io_input_payload_delay_13_stateElements_9 <= io_input_payload_delay_12_stateElements_9;
    io_input_payload_delay_13_stateElements_10 <= io_input_payload_delay_12_stateElements_10;
    io_input_payload_delay_13_stateElement <= io_input_payload_delay_12_stateElement;
    io_input_payload_delay_14_isFull <= io_input_payload_delay_13_isFull;
    io_input_payload_delay_14_fullRound <= io_input_payload_delay_13_fullRound;
    io_input_payload_delay_14_partialRound <= io_input_payload_delay_13_partialRound;
    io_input_payload_delay_14_stateIndex <= io_input_payload_delay_13_stateIndex;
    io_input_payload_delay_14_stateSize <= io_input_payload_delay_13_stateSize;
    io_input_payload_delay_14_stateID <= io_input_payload_delay_13_stateID;
    io_input_payload_delay_14_stateElements_0 <= io_input_payload_delay_13_stateElements_0;
    io_input_payload_delay_14_stateElements_1 <= io_input_payload_delay_13_stateElements_1;
    io_input_payload_delay_14_stateElements_2 <= io_input_payload_delay_13_stateElements_2;
    io_input_payload_delay_14_stateElements_3 <= io_input_payload_delay_13_stateElements_3;
    io_input_payload_delay_14_stateElements_4 <= io_input_payload_delay_13_stateElements_4;
    io_input_payload_delay_14_stateElements_5 <= io_input_payload_delay_13_stateElements_5;
    io_input_payload_delay_14_stateElements_6 <= io_input_payload_delay_13_stateElements_6;
    io_input_payload_delay_14_stateElements_7 <= io_input_payload_delay_13_stateElements_7;
    io_input_payload_delay_14_stateElements_8 <= io_input_payload_delay_13_stateElements_8;
    io_input_payload_delay_14_stateElements_9 <= io_input_payload_delay_13_stateElements_9;
    io_input_payload_delay_14_stateElements_10 <= io_input_payload_delay_13_stateElements_10;
    io_input_payload_delay_14_stateElement <= io_input_payload_delay_13_stateElement;
    io_input_payload_delay_15_isFull <= io_input_payload_delay_14_isFull;
    io_input_payload_delay_15_fullRound <= io_input_payload_delay_14_fullRound;
    io_input_payload_delay_15_partialRound <= io_input_payload_delay_14_partialRound;
    io_input_payload_delay_15_stateIndex <= io_input_payload_delay_14_stateIndex;
    io_input_payload_delay_15_stateSize <= io_input_payload_delay_14_stateSize;
    io_input_payload_delay_15_stateID <= io_input_payload_delay_14_stateID;
    io_input_payload_delay_15_stateElements_0 <= io_input_payload_delay_14_stateElements_0;
    io_input_payload_delay_15_stateElements_1 <= io_input_payload_delay_14_stateElements_1;
    io_input_payload_delay_15_stateElements_2 <= io_input_payload_delay_14_stateElements_2;
    io_input_payload_delay_15_stateElements_3 <= io_input_payload_delay_14_stateElements_3;
    io_input_payload_delay_15_stateElements_4 <= io_input_payload_delay_14_stateElements_4;
    io_input_payload_delay_15_stateElements_5 <= io_input_payload_delay_14_stateElements_5;
    io_input_payload_delay_15_stateElements_6 <= io_input_payload_delay_14_stateElements_6;
    io_input_payload_delay_15_stateElements_7 <= io_input_payload_delay_14_stateElements_7;
    io_input_payload_delay_15_stateElements_8 <= io_input_payload_delay_14_stateElements_8;
    io_input_payload_delay_15_stateElements_9 <= io_input_payload_delay_14_stateElements_9;
    io_input_payload_delay_15_stateElements_10 <= io_input_payload_delay_14_stateElements_10;
    io_input_payload_delay_15_stateElement <= io_input_payload_delay_14_stateElement;
    io_input_payload_delay_16_isFull <= io_input_payload_delay_15_isFull;
    io_input_payload_delay_16_fullRound <= io_input_payload_delay_15_fullRound;
    io_input_payload_delay_16_partialRound <= io_input_payload_delay_15_partialRound;
    io_input_payload_delay_16_stateIndex <= io_input_payload_delay_15_stateIndex;
    io_input_payload_delay_16_stateSize <= io_input_payload_delay_15_stateSize;
    io_input_payload_delay_16_stateID <= io_input_payload_delay_15_stateID;
    io_input_payload_delay_16_stateElements_0 <= io_input_payload_delay_15_stateElements_0;
    io_input_payload_delay_16_stateElements_1 <= io_input_payload_delay_15_stateElements_1;
    io_input_payload_delay_16_stateElements_2 <= io_input_payload_delay_15_stateElements_2;
    io_input_payload_delay_16_stateElements_3 <= io_input_payload_delay_15_stateElements_3;
    io_input_payload_delay_16_stateElements_4 <= io_input_payload_delay_15_stateElements_4;
    io_input_payload_delay_16_stateElements_5 <= io_input_payload_delay_15_stateElements_5;
    io_input_payload_delay_16_stateElements_6 <= io_input_payload_delay_15_stateElements_6;
    io_input_payload_delay_16_stateElements_7 <= io_input_payload_delay_15_stateElements_7;
    io_input_payload_delay_16_stateElements_8 <= io_input_payload_delay_15_stateElements_8;
    io_input_payload_delay_16_stateElements_9 <= io_input_payload_delay_15_stateElements_9;
    io_input_payload_delay_16_stateElements_10 <= io_input_payload_delay_15_stateElements_10;
    io_input_payload_delay_16_stateElement <= io_input_payload_delay_15_stateElement;
    io_input_payload_delay_17_isFull <= io_input_payload_delay_16_isFull;
    io_input_payload_delay_17_fullRound <= io_input_payload_delay_16_fullRound;
    io_input_payload_delay_17_partialRound <= io_input_payload_delay_16_partialRound;
    io_input_payload_delay_17_stateIndex <= io_input_payload_delay_16_stateIndex;
    io_input_payload_delay_17_stateSize <= io_input_payload_delay_16_stateSize;
    io_input_payload_delay_17_stateID <= io_input_payload_delay_16_stateID;
    io_input_payload_delay_17_stateElements_0 <= io_input_payload_delay_16_stateElements_0;
    io_input_payload_delay_17_stateElements_1 <= io_input_payload_delay_16_stateElements_1;
    io_input_payload_delay_17_stateElements_2 <= io_input_payload_delay_16_stateElements_2;
    io_input_payload_delay_17_stateElements_3 <= io_input_payload_delay_16_stateElements_3;
    io_input_payload_delay_17_stateElements_4 <= io_input_payload_delay_16_stateElements_4;
    io_input_payload_delay_17_stateElements_5 <= io_input_payload_delay_16_stateElements_5;
    io_input_payload_delay_17_stateElements_6 <= io_input_payload_delay_16_stateElements_6;
    io_input_payload_delay_17_stateElements_7 <= io_input_payload_delay_16_stateElements_7;
    io_input_payload_delay_17_stateElements_8 <= io_input_payload_delay_16_stateElements_8;
    io_input_payload_delay_17_stateElements_9 <= io_input_payload_delay_16_stateElements_9;
    io_input_payload_delay_17_stateElements_10 <= io_input_payload_delay_16_stateElements_10;
    io_input_payload_delay_17_stateElement <= io_input_payload_delay_16_stateElement;
    io_input_payload_delay_18_isFull <= io_input_payload_delay_17_isFull;
    io_input_payload_delay_18_fullRound <= io_input_payload_delay_17_fullRound;
    io_input_payload_delay_18_partialRound <= io_input_payload_delay_17_partialRound;
    io_input_payload_delay_18_stateIndex <= io_input_payload_delay_17_stateIndex;
    io_input_payload_delay_18_stateSize <= io_input_payload_delay_17_stateSize;
    io_input_payload_delay_18_stateID <= io_input_payload_delay_17_stateID;
    io_input_payload_delay_18_stateElements_0 <= io_input_payload_delay_17_stateElements_0;
    io_input_payload_delay_18_stateElements_1 <= io_input_payload_delay_17_stateElements_1;
    io_input_payload_delay_18_stateElements_2 <= io_input_payload_delay_17_stateElements_2;
    io_input_payload_delay_18_stateElements_3 <= io_input_payload_delay_17_stateElements_3;
    io_input_payload_delay_18_stateElements_4 <= io_input_payload_delay_17_stateElements_4;
    io_input_payload_delay_18_stateElements_5 <= io_input_payload_delay_17_stateElements_5;
    io_input_payload_delay_18_stateElements_6 <= io_input_payload_delay_17_stateElements_6;
    io_input_payload_delay_18_stateElements_7 <= io_input_payload_delay_17_stateElements_7;
    io_input_payload_delay_18_stateElements_8 <= io_input_payload_delay_17_stateElements_8;
    io_input_payload_delay_18_stateElements_9 <= io_input_payload_delay_17_stateElements_9;
    io_input_payload_delay_18_stateElements_10 <= io_input_payload_delay_17_stateElements_10;
    io_input_payload_delay_18_stateElement <= io_input_payload_delay_17_stateElement;
    io_input_payload_delay_19_isFull <= io_input_payload_delay_18_isFull;
    io_input_payload_delay_19_fullRound <= io_input_payload_delay_18_fullRound;
    io_input_payload_delay_19_partialRound <= io_input_payload_delay_18_partialRound;
    io_input_payload_delay_19_stateIndex <= io_input_payload_delay_18_stateIndex;
    io_input_payload_delay_19_stateSize <= io_input_payload_delay_18_stateSize;
    io_input_payload_delay_19_stateID <= io_input_payload_delay_18_stateID;
    io_input_payload_delay_19_stateElements_0 <= io_input_payload_delay_18_stateElements_0;
    io_input_payload_delay_19_stateElements_1 <= io_input_payload_delay_18_stateElements_1;
    io_input_payload_delay_19_stateElements_2 <= io_input_payload_delay_18_stateElements_2;
    io_input_payload_delay_19_stateElements_3 <= io_input_payload_delay_18_stateElements_3;
    io_input_payload_delay_19_stateElements_4 <= io_input_payload_delay_18_stateElements_4;
    io_input_payload_delay_19_stateElements_5 <= io_input_payload_delay_18_stateElements_5;
    io_input_payload_delay_19_stateElements_6 <= io_input_payload_delay_18_stateElements_6;
    io_input_payload_delay_19_stateElements_7 <= io_input_payload_delay_18_stateElements_7;
    io_input_payload_delay_19_stateElements_8 <= io_input_payload_delay_18_stateElements_8;
    io_input_payload_delay_19_stateElements_9 <= io_input_payload_delay_18_stateElements_9;
    io_input_payload_delay_19_stateElements_10 <= io_input_payload_delay_18_stateElements_10;
    io_input_payload_delay_19_stateElement <= io_input_payload_delay_18_stateElement;
    io_input_payload_delay_20_isFull <= io_input_payload_delay_19_isFull;
    io_input_payload_delay_20_fullRound <= io_input_payload_delay_19_fullRound;
    io_input_payload_delay_20_partialRound <= io_input_payload_delay_19_partialRound;
    io_input_payload_delay_20_stateIndex <= io_input_payload_delay_19_stateIndex;
    io_input_payload_delay_20_stateSize <= io_input_payload_delay_19_stateSize;
    io_input_payload_delay_20_stateID <= io_input_payload_delay_19_stateID;
    io_input_payload_delay_20_stateElements_0 <= io_input_payload_delay_19_stateElements_0;
    io_input_payload_delay_20_stateElements_1 <= io_input_payload_delay_19_stateElements_1;
    io_input_payload_delay_20_stateElements_2 <= io_input_payload_delay_19_stateElements_2;
    io_input_payload_delay_20_stateElements_3 <= io_input_payload_delay_19_stateElements_3;
    io_input_payload_delay_20_stateElements_4 <= io_input_payload_delay_19_stateElements_4;
    io_input_payload_delay_20_stateElements_5 <= io_input_payload_delay_19_stateElements_5;
    io_input_payload_delay_20_stateElements_6 <= io_input_payload_delay_19_stateElements_6;
    io_input_payload_delay_20_stateElements_7 <= io_input_payload_delay_19_stateElements_7;
    io_input_payload_delay_20_stateElements_8 <= io_input_payload_delay_19_stateElements_8;
    io_input_payload_delay_20_stateElements_9 <= io_input_payload_delay_19_stateElements_9;
    io_input_payload_delay_20_stateElements_10 <= io_input_payload_delay_19_stateElements_10;
    io_input_payload_delay_20_stateElement <= io_input_payload_delay_19_stateElement;
    io_input_payload_delay_21_isFull <= io_input_payload_delay_20_isFull;
    io_input_payload_delay_21_fullRound <= io_input_payload_delay_20_fullRound;
    io_input_payload_delay_21_partialRound <= io_input_payload_delay_20_partialRound;
    io_input_payload_delay_21_stateIndex <= io_input_payload_delay_20_stateIndex;
    io_input_payload_delay_21_stateSize <= io_input_payload_delay_20_stateSize;
    io_input_payload_delay_21_stateID <= io_input_payload_delay_20_stateID;
    io_input_payload_delay_21_stateElements_0 <= io_input_payload_delay_20_stateElements_0;
    io_input_payload_delay_21_stateElements_1 <= io_input_payload_delay_20_stateElements_1;
    io_input_payload_delay_21_stateElements_2 <= io_input_payload_delay_20_stateElements_2;
    io_input_payload_delay_21_stateElements_3 <= io_input_payload_delay_20_stateElements_3;
    io_input_payload_delay_21_stateElements_4 <= io_input_payload_delay_20_stateElements_4;
    io_input_payload_delay_21_stateElements_5 <= io_input_payload_delay_20_stateElements_5;
    io_input_payload_delay_21_stateElements_6 <= io_input_payload_delay_20_stateElements_6;
    io_input_payload_delay_21_stateElements_7 <= io_input_payload_delay_20_stateElements_7;
    io_input_payload_delay_21_stateElements_8 <= io_input_payload_delay_20_stateElements_8;
    io_input_payload_delay_21_stateElements_9 <= io_input_payload_delay_20_stateElements_9;
    io_input_payload_delay_21_stateElements_10 <= io_input_payload_delay_20_stateElements_10;
    io_input_payload_delay_21_stateElement <= io_input_payload_delay_20_stateElement;
    io_input_payload_delay_22_isFull <= io_input_payload_delay_21_isFull;
    io_input_payload_delay_22_fullRound <= io_input_payload_delay_21_fullRound;
    io_input_payload_delay_22_partialRound <= io_input_payload_delay_21_partialRound;
    io_input_payload_delay_22_stateIndex <= io_input_payload_delay_21_stateIndex;
    io_input_payload_delay_22_stateSize <= io_input_payload_delay_21_stateSize;
    io_input_payload_delay_22_stateID <= io_input_payload_delay_21_stateID;
    io_input_payload_delay_22_stateElements_0 <= io_input_payload_delay_21_stateElements_0;
    io_input_payload_delay_22_stateElements_1 <= io_input_payload_delay_21_stateElements_1;
    io_input_payload_delay_22_stateElements_2 <= io_input_payload_delay_21_stateElements_2;
    io_input_payload_delay_22_stateElements_3 <= io_input_payload_delay_21_stateElements_3;
    io_input_payload_delay_22_stateElements_4 <= io_input_payload_delay_21_stateElements_4;
    io_input_payload_delay_22_stateElements_5 <= io_input_payload_delay_21_stateElements_5;
    io_input_payload_delay_22_stateElements_6 <= io_input_payload_delay_21_stateElements_6;
    io_input_payload_delay_22_stateElements_7 <= io_input_payload_delay_21_stateElements_7;
    io_input_payload_delay_22_stateElements_8 <= io_input_payload_delay_21_stateElements_8;
    io_input_payload_delay_22_stateElements_9 <= io_input_payload_delay_21_stateElements_9;
    io_input_payload_delay_22_stateElements_10 <= io_input_payload_delay_21_stateElements_10;
    io_input_payload_delay_22_stateElement <= io_input_payload_delay_21_stateElement;
    io_input_payload_delay_23_isFull <= io_input_payload_delay_22_isFull;
    io_input_payload_delay_23_fullRound <= io_input_payload_delay_22_fullRound;
    io_input_payload_delay_23_partialRound <= io_input_payload_delay_22_partialRound;
    io_input_payload_delay_23_stateIndex <= io_input_payload_delay_22_stateIndex;
    io_input_payload_delay_23_stateSize <= io_input_payload_delay_22_stateSize;
    io_input_payload_delay_23_stateID <= io_input_payload_delay_22_stateID;
    io_input_payload_delay_23_stateElements_0 <= io_input_payload_delay_22_stateElements_0;
    io_input_payload_delay_23_stateElements_1 <= io_input_payload_delay_22_stateElements_1;
    io_input_payload_delay_23_stateElements_2 <= io_input_payload_delay_22_stateElements_2;
    io_input_payload_delay_23_stateElements_3 <= io_input_payload_delay_22_stateElements_3;
    io_input_payload_delay_23_stateElements_4 <= io_input_payload_delay_22_stateElements_4;
    io_input_payload_delay_23_stateElements_5 <= io_input_payload_delay_22_stateElements_5;
    io_input_payload_delay_23_stateElements_6 <= io_input_payload_delay_22_stateElements_6;
    io_input_payload_delay_23_stateElements_7 <= io_input_payload_delay_22_stateElements_7;
    io_input_payload_delay_23_stateElements_8 <= io_input_payload_delay_22_stateElements_8;
    io_input_payload_delay_23_stateElements_9 <= io_input_payload_delay_22_stateElements_9;
    io_input_payload_delay_23_stateElements_10 <= io_input_payload_delay_22_stateElements_10;
    io_input_payload_delay_23_stateElement <= io_input_payload_delay_22_stateElement;
    io_input_payload_delay_24_isFull <= io_input_payload_delay_23_isFull;
    io_input_payload_delay_24_fullRound <= io_input_payload_delay_23_fullRound;
    io_input_payload_delay_24_partialRound <= io_input_payload_delay_23_partialRound;
    io_input_payload_delay_24_stateIndex <= io_input_payload_delay_23_stateIndex;
    io_input_payload_delay_24_stateSize <= io_input_payload_delay_23_stateSize;
    io_input_payload_delay_24_stateID <= io_input_payload_delay_23_stateID;
    io_input_payload_delay_24_stateElements_0 <= io_input_payload_delay_23_stateElements_0;
    io_input_payload_delay_24_stateElements_1 <= io_input_payload_delay_23_stateElements_1;
    io_input_payload_delay_24_stateElements_2 <= io_input_payload_delay_23_stateElements_2;
    io_input_payload_delay_24_stateElements_3 <= io_input_payload_delay_23_stateElements_3;
    io_input_payload_delay_24_stateElements_4 <= io_input_payload_delay_23_stateElements_4;
    io_input_payload_delay_24_stateElements_5 <= io_input_payload_delay_23_stateElements_5;
    io_input_payload_delay_24_stateElements_6 <= io_input_payload_delay_23_stateElements_6;
    io_input_payload_delay_24_stateElements_7 <= io_input_payload_delay_23_stateElements_7;
    io_input_payload_delay_24_stateElements_8 <= io_input_payload_delay_23_stateElements_8;
    io_input_payload_delay_24_stateElements_9 <= io_input_payload_delay_23_stateElements_9;
    io_input_payload_delay_24_stateElements_10 <= io_input_payload_delay_23_stateElements_10;
    io_input_payload_delay_24_stateElement <= io_input_payload_delay_23_stateElement;
    io_input_payload_delay_25_isFull <= io_input_payload_delay_24_isFull;
    io_input_payload_delay_25_fullRound <= io_input_payload_delay_24_fullRound;
    io_input_payload_delay_25_partialRound <= io_input_payload_delay_24_partialRound;
    io_input_payload_delay_25_stateIndex <= io_input_payload_delay_24_stateIndex;
    io_input_payload_delay_25_stateSize <= io_input_payload_delay_24_stateSize;
    io_input_payload_delay_25_stateID <= io_input_payload_delay_24_stateID;
    io_input_payload_delay_25_stateElements_0 <= io_input_payload_delay_24_stateElements_0;
    io_input_payload_delay_25_stateElements_1 <= io_input_payload_delay_24_stateElements_1;
    io_input_payload_delay_25_stateElements_2 <= io_input_payload_delay_24_stateElements_2;
    io_input_payload_delay_25_stateElements_3 <= io_input_payload_delay_24_stateElements_3;
    io_input_payload_delay_25_stateElements_4 <= io_input_payload_delay_24_stateElements_4;
    io_input_payload_delay_25_stateElements_5 <= io_input_payload_delay_24_stateElements_5;
    io_input_payload_delay_25_stateElements_6 <= io_input_payload_delay_24_stateElements_6;
    io_input_payload_delay_25_stateElements_7 <= io_input_payload_delay_24_stateElements_7;
    io_input_payload_delay_25_stateElements_8 <= io_input_payload_delay_24_stateElements_8;
    io_input_payload_delay_25_stateElements_9 <= io_input_payload_delay_24_stateElements_9;
    io_input_payload_delay_25_stateElements_10 <= io_input_payload_delay_24_stateElements_10;
    io_input_payload_delay_25_stateElement <= io_input_payload_delay_24_stateElement;
    io_input_payload_delay_26_isFull <= io_input_payload_delay_25_isFull;
    io_input_payload_delay_26_fullRound <= io_input_payload_delay_25_fullRound;
    io_input_payload_delay_26_partialRound <= io_input_payload_delay_25_partialRound;
    io_input_payload_delay_26_stateIndex <= io_input_payload_delay_25_stateIndex;
    io_input_payload_delay_26_stateSize <= io_input_payload_delay_25_stateSize;
    io_input_payload_delay_26_stateID <= io_input_payload_delay_25_stateID;
    io_input_payload_delay_26_stateElements_0 <= io_input_payload_delay_25_stateElements_0;
    io_input_payload_delay_26_stateElements_1 <= io_input_payload_delay_25_stateElements_1;
    io_input_payload_delay_26_stateElements_2 <= io_input_payload_delay_25_stateElements_2;
    io_input_payload_delay_26_stateElements_3 <= io_input_payload_delay_25_stateElements_3;
    io_input_payload_delay_26_stateElements_4 <= io_input_payload_delay_25_stateElements_4;
    io_input_payload_delay_26_stateElements_5 <= io_input_payload_delay_25_stateElements_5;
    io_input_payload_delay_26_stateElements_6 <= io_input_payload_delay_25_stateElements_6;
    io_input_payload_delay_26_stateElements_7 <= io_input_payload_delay_25_stateElements_7;
    io_input_payload_delay_26_stateElements_8 <= io_input_payload_delay_25_stateElements_8;
    io_input_payload_delay_26_stateElements_9 <= io_input_payload_delay_25_stateElements_9;
    io_input_payload_delay_26_stateElements_10 <= io_input_payload_delay_25_stateElements_10;
    io_input_payload_delay_26_stateElement <= io_input_payload_delay_25_stateElement;
    io_input_payload_delay_27_isFull <= io_input_payload_delay_26_isFull;
    io_input_payload_delay_27_fullRound <= io_input_payload_delay_26_fullRound;
    io_input_payload_delay_27_partialRound <= io_input_payload_delay_26_partialRound;
    io_input_payload_delay_27_stateIndex <= io_input_payload_delay_26_stateIndex;
    io_input_payload_delay_27_stateSize <= io_input_payload_delay_26_stateSize;
    io_input_payload_delay_27_stateID <= io_input_payload_delay_26_stateID;
    io_input_payload_delay_27_stateElements_0 <= io_input_payload_delay_26_stateElements_0;
    io_input_payload_delay_27_stateElements_1 <= io_input_payload_delay_26_stateElements_1;
    io_input_payload_delay_27_stateElements_2 <= io_input_payload_delay_26_stateElements_2;
    io_input_payload_delay_27_stateElements_3 <= io_input_payload_delay_26_stateElements_3;
    io_input_payload_delay_27_stateElements_4 <= io_input_payload_delay_26_stateElements_4;
    io_input_payload_delay_27_stateElements_5 <= io_input_payload_delay_26_stateElements_5;
    io_input_payload_delay_27_stateElements_6 <= io_input_payload_delay_26_stateElements_6;
    io_input_payload_delay_27_stateElements_7 <= io_input_payload_delay_26_stateElements_7;
    io_input_payload_delay_27_stateElements_8 <= io_input_payload_delay_26_stateElements_8;
    io_input_payload_delay_27_stateElements_9 <= io_input_payload_delay_26_stateElements_9;
    io_input_payload_delay_27_stateElements_10 <= io_input_payload_delay_26_stateElements_10;
    io_input_payload_delay_27_stateElement <= io_input_payload_delay_26_stateElement;
    io_input_payload_delay_28_isFull <= io_input_payload_delay_27_isFull;
    io_input_payload_delay_28_fullRound <= io_input_payload_delay_27_fullRound;
    io_input_payload_delay_28_partialRound <= io_input_payload_delay_27_partialRound;
    io_input_payload_delay_28_stateIndex <= io_input_payload_delay_27_stateIndex;
    io_input_payload_delay_28_stateSize <= io_input_payload_delay_27_stateSize;
    io_input_payload_delay_28_stateID <= io_input_payload_delay_27_stateID;
    io_input_payload_delay_28_stateElements_0 <= io_input_payload_delay_27_stateElements_0;
    io_input_payload_delay_28_stateElements_1 <= io_input_payload_delay_27_stateElements_1;
    io_input_payload_delay_28_stateElements_2 <= io_input_payload_delay_27_stateElements_2;
    io_input_payload_delay_28_stateElements_3 <= io_input_payload_delay_27_stateElements_3;
    io_input_payload_delay_28_stateElements_4 <= io_input_payload_delay_27_stateElements_4;
    io_input_payload_delay_28_stateElements_5 <= io_input_payload_delay_27_stateElements_5;
    io_input_payload_delay_28_stateElements_6 <= io_input_payload_delay_27_stateElements_6;
    io_input_payload_delay_28_stateElements_7 <= io_input_payload_delay_27_stateElements_7;
    io_input_payload_delay_28_stateElements_8 <= io_input_payload_delay_27_stateElements_8;
    io_input_payload_delay_28_stateElements_9 <= io_input_payload_delay_27_stateElements_9;
    io_input_payload_delay_28_stateElements_10 <= io_input_payload_delay_27_stateElements_10;
    io_input_payload_delay_28_stateElement <= io_input_payload_delay_27_stateElement;
    io_input_payload_delay_29_isFull <= io_input_payload_delay_28_isFull;
    io_input_payload_delay_29_fullRound <= io_input_payload_delay_28_fullRound;
    io_input_payload_delay_29_partialRound <= io_input_payload_delay_28_partialRound;
    io_input_payload_delay_29_stateIndex <= io_input_payload_delay_28_stateIndex;
    io_input_payload_delay_29_stateSize <= io_input_payload_delay_28_stateSize;
    io_input_payload_delay_29_stateID <= io_input_payload_delay_28_stateID;
    io_input_payload_delay_29_stateElements_0 <= io_input_payload_delay_28_stateElements_0;
    io_input_payload_delay_29_stateElements_1 <= io_input_payload_delay_28_stateElements_1;
    io_input_payload_delay_29_stateElements_2 <= io_input_payload_delay_28_stateElements_2;
    io_input_payload_delay_29_stateElements_3 <= io_input_payload_delay_28_stateElements_3;
    io_input_payload_delay_29_stateElements_4 <= io_input_payload_delay_28_stateElements_4;
    io_input_payload_delay_29_stateElements_5 <= io_input_payload_delay_28_stateElements_5;
    io_input_payload_delay_29_stateElements_6 <= io_input_payload_delay_28_stateElements_6;
    io_input_payload_delay_29_stateElements_7 <= io_input_payload_delay_28_stateElements_7;
    io_input_payload_delay_29_stateElements_8 <= io_input_payload_delay_28_stateElements_8;
    io_input_payload_delay_29_stateElements_9 <= io_input_payload_delay_28_stateElements_9;
    io_input_payload_delay_29_stateElements_10 <= io_input_payload_delay_28_stateElements_10;
    io_input_payload_delay_29_stateElement <= io_input_payload_delay_28_stateElement;
    io_input_payload_delay_30_isFull <= io_input_payload_delay_29_isFull;
    io_input_payload_delay_30_fullRound <= io_input_payload_delay_29_fullRound;
    io_input_payload_delay_30_partialRound <= io_input_payload_delay_29_partialRound;
    io_input_payload_delay_30_stateIndex <= io_input_payload_delay_29_stateIndex;
    io_input_payload_delay_30_stateSize <= io_input_payload_delay_29_stateSize;
    io_input_payload_delay_30_stateID <= io_input_payload_delay_29_stateID;
    io_input_payload_delay_30_stateElements_0 <= io_input_payload_delay_29_stateElements_0;
    io_input_payload_delay_30_stateElements_1 <= io_input_payload_delay_29_stateElements_1;
    io_input_payload_delay_30_stateElements_2 <= io_input_payload_delay_29_stateElements_2;
    io_input_payload_delay_30_stateElements_3 <= io_input_payload_delay_29_stateElements_3;
    io_input_payload_delay_30_stateElements_4 <= io_input_payload_delay_29_stateElements_4;
    io_input_payload_delay_30_stateElements_5 <= io_input_payload_delay_29_stateElements_5;
    io_input_payload_delay_30_stateElements_6 <= io_input_payload_delay_29_stateElements_6;
    io_input_payload_delay_30_stateElements_7 <= io_input_payload_delay_29_stateElements_7;
    io_input_payload_delay_30_stateElements_8 <= io_input_payload_delay_29_stateElements_8;
    io_input_payload_delay_30_stateElements_9 <= io_input_payload_delay_29_stateElements_9;
    io_input_payload_delay_30_stateElements_10 <= io_input_payload_delay_29_stateElements_10;
    io_input_payload_delay_30_stateElement <= io_input_payload_delay_29_stateElement;
    io_input_payload_delay_31_isFull <= io_input_payload_delay_30_isFull;
    io_input_payload_delay_31_fullRound <= io_input_payload_delay_30_fullRound;
    io_input_payload_delay_31_partialRound <= io_input_payload_delay_30_partialRound;
    io_input_payload_delay_31_stateIndex <= io_input_payload_delay_30_stateIndex;
    io_input_payload_delay_31_stateSize <= io_input_payload_delay_30_stateSize;
    io_input_payload_delay_31_stateID <= io_input_payload_delay_30_stateID;
    io_input_payload_delay_31_stateElements_0 <= io_input_payload_delay_30_stateElements_0;
    io_input_payload_delay_31_stateElements_1 <= io_input_payload_delay_30_stateElements_1;
    io_input_payload_delay_31_stateElements_2 <= io_input_payload_delay_30_stateElements_2;
    io_input_payload_delay_31_stateElements_3 <= io_input_payload_delay_30_stateElements_3;
    io_input_payload_delay_31_stateElements_4 <= io_input_payload_delay_30_stateElements_4;
    io_input_payload_delay_31_stateElements_5 <= io_input_payload_delay_30_stateElements_5;
    io_input_payload_delay_31_stateElements_6 <= io_input_payload_delay_30_stateElements_6;
    io_input_payload_delay_31_stateElements_7 <= io_input_payload_delay_30_stateElements_7;
    io_input_payload_delay_31_stateElements_8 <= io_input_payload_delay_30_stateElements_8;
    io_input_payload_delay_31_stateElements_9 <= io_input_payload_delay_30_stateElements_9;
    io_input_payload_delay_31_stateElements_10 <= io_input_payload_delay_30_stateElements_10;
    io_input_payload_delay_31_stateElement <= io_input_payload_delay_30_stateElement;
    io_input_payload_delay_32_isFull <= io_input_payload_delay_31_isFull;
    io_input_payload_delay_32_fullRound <= io_input_payload_delay_31_fullRound;
    io_input_payload_delay_32_partialRound <= io_input_payload_delay_31_partialRound;
    io_input_payload_delay_32_stateIndex <= io_input_payload_delay_31_stateIndex;
    io_input_payload_delay_32_stateSize <= io_input_payload_delay_31_stateSize;
    io_input_payload_delay_32_stateID <= io_input_payload_delay_31_stateID;
    io_input_payload_delay_32_stateElements_0 <= io_input_payload_delay_31_stateElements_0;
    io_input_payload_delay_32_stateElements_1 <= io_input_payload_delay_31_stateElements_1;
    io_input_payload_delay_32_stateElements_2 <= io_input_payload_delay_31_stateElements_2;
    io_input_payload_delay_32_stateElements_3 <= io_input_payload_delay_31_stateElements_3;
    io_input_payload_delay_32_stateElements_4 <= io_input_payload_delay_31_stateElements_4;
    io_input_payload_delay_32_stateElements_5 <= io_input_payload_delay_31_stateElements_5;
    io_input_payload_delay_32_stateElements_6 <= io_input_payload_delay_31_stateElements_6;
    io_input_payload_delay_32_stateElements_7 <= io_input_payload_delay_31_stateElements_7;
    io_input_payload_delay_32_stateElements_8 <= io_input_payload_delay_31_stateElements_8;
    io_input_payload_delay_32_stateElements_9 <= io_input_payload_delay_31_stateElements_9;
    io_input_payload_delay_32_stateElements_10 <= io_input_payload_delay_31_stateElements_10;
    io_input_payload_delay_32_stateElement <= io_input_payload_delay_31_stateElement;
    io_input_payload_delay_33_isFull <= io_input_payload_delay_32_isFull;
    io_input_payload_delay_33_fullRound <= io_input_payload_delay_32_fullRound;
    io_input_payload_delay_33_partialRound <= io_input_payload_delay_32_partialRound;
    io_input_payload_delay_33_stateIndex <= io_input_payload_delay_32_stateIndex;
    io_input_payload_delay_33_stateSize <= io_input_payload_delay_32_stateSize;
    io_input_payload_delay_33_stateID <= io_input_payload_delay_32_stateID;
    io_input_payload_delay_33_stateElements_0 <= io_input_payload_delay_32_stateElements_0;
    io_input_payload_delay_33_stateElements_1 <= io_input_payload_delay_32_stateElements_1;
    io_input_payload_delay_33_stateElements_2 <= io_input_payload_delay_32_stateElements_2;
    io_input_payload_delay_33_stateElements_3 <= io_input_payload_delay_32_stateElements_3;
    io_input_payload_delay_33_stateElements_4 <= io_input_payload_delay_32_stateElements_4;
    io_input_payload_delay_33_stateElements_5 <= io_input_payload_delay_32_stateElements_5;
    io_input_payload_delay_33_stateElements_6 <= io_input_payload_delay_32_stateElements_6;
    io_input_payload_delay_33_stateElements_7 <= io_input_payload_delay_32_stateElements_7;
    io_input_payload_delay_33_stateElements_8 <= io_input_payload_delay_32_stateElements_8;
    io_input_payload_delay_33_stateElements_9 <= io_input_payload_delay_32_stateElements_9;
    io_input_payload_delay_33_stateElements_10 <= io_input_payload_delay_32_stateElements_10;
    io_input_payload_delay_33_stateElement <= io_input_payload_delay_32_stateElement;
    io_input_payload_delay_34_isFull <= io_input_payload_delay_33_isFull;
    io_input_payload_delay_34_fullRound <= io_input_payload_delay_33_fullRound;
    io_input_payload_delay_34_partialRound <= io_input_payload_delay_33_partialRound;
    io_input_payload_delay_34_stateIndex <= io_input_payload_delay_33_stateIndex;
    io_input_payload_delay_34_stateSize <= io_input_payload_delay_33_stateSize;
    io_input_payload_delay_34_stateID <= io_input_payload_delay_33_stateID;
    io_input_payload_delay_34_stateElements_0 <= io_input_payload_delay_33_stateElements_0;
    io_input_payload_delay_34_stateElements_1 <= io_input_payload_delay_33_stateElements_1;
    io_input_payload_delay_34_stateElements_2 <= io_input_payload_delay_33_stateElements_2;
    io_input_payload_delay_34_stateElements_3 <= io_input_payload_delay_33_stateElements_3;
    io_input_payload_delay_34_stateElements_4 <= io_input_payload_delay_33_stateElements_4;
    io_input_payload_delay_34_stateElements_5 <= io_input_payload_delay_33_stateElements_5;
    io_input_payload_delay_34_stateElements_6 <= io_input_payload_delay_33_stateElements_6;
    io_input_payload_delay_34_stateElements_7 <= io_input_payload_delay_33_stateElements_7;
    io_input_payload_delay_34_stateElements_8 <= io_input_payload_delay_33_stateElements_8;
    io_input_payload_delay_34_stateElements_9 <= io_input_payload_delay_33_stateElements_9;
    io_input_payload_delay_34_stateElements_10 <= io_input_payload_delay_33_stateElements_10;
    io_input_payload_delay_34_stateElement <= io_input_payload_delay_33_stateElement;
    io_input_payload_delay_35_isFull <= io_input_payload_delay_34_isFull;
    io_input_payload_delay_35_fullRound <= io_input_payload_delay_34_fullRound;
    io_input_payload_delay_35_partialRound <= io_input_payload_delay_34_partialRound;
    io_input_payload_delay_35_stateIndex <= io_input_payload_delay_34_stateIndex;
    io_input_payload_delay_35_stateSize <= io_input_payload_delay_34_stateSize;
    io_input_payload_delay_35_stateID <= io_input_payload_delay_34_stateID;
    io_input_payload_delay_35_stateElements_0 <= io_input_payload_delay_34_stateElements_0;
    io_input_payload_delay_35_stateElements_1 <= io_input_payload_delay_34_stateElements_1;
    io_input_payload_delay_35_stateElements_2 <= io_input_payload_delay_34_stateElements_2;
    io_input_payload_delay_35_stateElements_3 <= io_input_payload_delay_34_stateElements_3;
    io_input_payload_delay_35_stateElements_4 <= io_input_payload_delay_34_stateElements_4;
    io_input_payload_delay_35_stateElements_5 <= io_input_payload_delay_34_stateElements_5;
    io_input_payload_delay_35_stateElements_6 <= io_input_payload_delay_34_stateElements_6;
    io_input_payload_delay_35_stateElements_7 <= io_input_payload_delay_34_stateElements_7;
    io_input_payload_delay_35_stateElements_8 <= io_input_payload_delay_34_stateElements_8;
    io_input_payload_delay_35_stateElements_9 <= io_input_payload_delay_34_stateElements_9;
    io_input_payload_delay_35_stateElements_10 <= io_input_payload_delay_34_stateElements_10;
    io_input_payload_delay_35_stateElement <= io_input_payload_delay_34_stateElement;
    io_input_payload_delay_36_isFull <= io_input_payload_delay_35_isFull;
    io_input_payload_delay_36_fullRound <= io_input_payload_delay_35_fullRound;
    io_input_payload_delay_36_partialRound <= io_input_payload_delay_35_partialRound;
    io_input_payload_delay_36_stateIndex <= io_input_payload_delay_35_stateIndex;
    io_input_payload_delay_36_stateSize <= io_input_payload_delay_35_stateSize;
    io_input_payload_delay_36_stateID <= io_input_payload_delay_35_stateID;
    io_input_payload_delay_36_stateElements_0 <= io_input_payload_delay_35_stateElements_0;
    io_input_payload_delay_36_stateElements_1 <= io_input_payload_delay_35_stateElements_1;
    io_input_payload_delay_36_stateElements_2 <= io_input_payload_delay_35_stateElements_2;
    io_input_payload_delay_36_stateElements_3 <= io_input_payload_delay_35_stateElements_3;
    io_input_payload_delay_36_stateElements_4 <= io_input_payload_delay_35_stateElements_4;
    io_input_payload_delay_36_stateElements_5 <= io_input_payload_delay_35_stateElements_5;
    io_input_payload_delay_36_stateElements_6 <= io_input_payload_delay_35_stateElements_6;
    io_input_payload_delay_36_stateElements_7 <= io_input_payload_delay_35_stateElements_7;
    io_input_payload_delay_36_stateElements_8 <= io_input_payload_delay_35_stateElements_8;
    io_input_payload_delay_36_stateElements_9 <= io_input_payload_delay_35_stateElements_9;
    io_input_payload_delay_36_stateElements_10 <= io_input_payload_delay_35_stateElements_10;
    io_input_payload_delay_36_stateElement <= io_input_payload_delay_35_stateElement;
    io_input_payload_delay_37_isFull <= io_input_payload_delay_36_isFull;
    io_input_payload_delay_37_fullRound <= io_input_payload_delay_36_fullRound;
    io_input_payload_delay_37_partialRound <= io_input_payload_delay_36_partialRound;
    io_input_payload_delay_37_stateIndex <= io_input_payload_delay_36_stateIndex;
    io_input_payload_delay_37_stateSize <= io_input_payload_delay_36_stateSize;
    io_input_payload_delay_37_stateID <= io_input_payload_delay_36_stateID;
    io_input_payload_delay_37_stateElements_0 <= io_input_payload_delay_36_stateElements_0;
    io_input_payload_delay_37_stateElements_1 <= io_input_payload_delay_36_stateElements_1;
    io_input_payload_delay_37_stateElements_2 <= io_input_payload_delay_36_stateElements_2;
    io_input_payload_delay_37_stateElements_3 <= io_input_payload_delay_36_stateElements_3;
    io_input_payload_delay_37_stateElements_4 <= io_input_payload_delay_36_stateElements_4;
    io_input_payload_delay_37_stateElements_5 <= io_input_payload_delay_36_stateElements_5;
    io_input_payload_delay_37_stateElements_6 <= io_input_payload_delay_36_stateElements_6;
    io_input_payload_delay_37_stateElements_7 <= io_input_payload_delay_36_stateElements_7;
    io_input_payload_delay_37_stateElements_8 <= io_input_payload_delay_36_stateElements_8;
    io_input_payload_delay_37_stateElements_9 <= io_input_payload_delay_36_stateElements_9;
    io_input_payload_delay_37_stateElements_10 <= io_input_payload_delay_36_stateElements_10;
    io_input_payload_delay_37_stateElement <= io_input_payload_delay_36_stateElement;
    io_input_payload_delay_38_isFull <= io_input_payload_delay_37_isFull;
    io_input_payload_delay_38_fullRound <= io_input_payload_delay_37_fullRound;
    io_input_payload_delay_38_partialRound <= io_input_payload_delay_37_partialRound;
    io_input_payload_delay_38_stateIndex <= io_input_payload_delay_37_stateIndex;
    io_input_payload_delay_38_stateSize <= io_input_payload_delay_37_stateSize;
    io_input_payload_delay_38_stateID <= io_input_payload_delay_37_stateID;
    io_input_payload_delay_38_stateElements_0 <= io_input_payload_delay_37_stateElements_0;
    io_input_payload_delay_38_stateElements_1 <= io_input_payload_delay_37_stateElements_1;
    io_input_payload_delay_38_stateElements_2 <= io_input_payload_delay_37_stateElements_2;
    io_input_payload_delay_38_stateElements_3 <= io_input_payload_delay_37_stateElements_3;
    io_input_payload_delay_38_stateElements_4 <= io_input_payload_delay_37_stateElements_4;
    io_input_payload_delay_38_stateElements_5 <= io_input_payload_delay_37_stateElements_5;
    io_input_payload_delay_38_stateElements_6 <= io_input_payload_delay_37_stateElements_6;
    io_input_payload_delay_38_stateElements_7 <= io_input_payload_delay_37_stateElements_7;
    io_input_payload_delay_38_stateElements_8 <= io_input_payload_delay_37_stateElements_8;
    io_input_payload_delay_38_stateElements_9 <= io_input_payload_delay_37_stateElements_9;
    io_input_payload_delay_38_stateElements_10 <= io_input_payload_delay_37_stateElements_10;
    io_input_payload_delay_38_stateElement <= io_input_payload_delay_37_stateElement;
    io_input_payload_delay_39_isFull <= io_input_payload_delay_38_isFull;
    io_input_payload_delay_39_fullRound <= io_input_payload_delay_38_fullRound;
    io_input_payload_delay_39_partialRound <= io_input_payload_delay_38_partialRound;
    io_input_payload_delay_39_stateIndex <= io_input_payload_delay_38_stateIndex;
    io_input_payload_delay_39_stateSize <= io_input_payload_delay_38_stateSize;
    io_input_payload_delay_39_stateID <= io_input_payload_delay_38_stateID;
    io_input_payload_delay_39_stateElements_0 <= io_input_payload_delay_38_stateElements_0;
    io_input_payload_delay_39_stateElements_1 <= io_input_payload_delay_38_stateElements_1;
    io_input_payload_delay_39_stateElements_2 <= io_input_payload_delay_38_stateElements_2;
    io_input_payload_delay_39_stateElements_3 <= io_input_payload_delay_38_stateElements_3;
    io_input_payload_delay_39_stateElements_4 <= io_input_payload_delay_38_stateElements_4;
    io_input_payload_delay_39_stateElements_5 <= io_input_payload_delay_38_stateElements_5;
    io_input_payload_delay_39_stateElements_6 <= io_input_payload_delay_38_stateElements_6;
    io_input_payload_delay_39_stateElements_7 <= io_input_payload_delay_38_stateElements_7;
    io_input_payload_delay_39_stateElements_8 <= io_input_payload_delay_38_stateElements_8;
    io_input_payload_delay_39_stateElements_9 <= io_input_payload_delay_38_stateElements_9;
    io_input_payload_delay_39_stateElements_10 <= io_input_payload_delay_38_stateElements_10;
    io_input_payload_delay_39_stateElement <= io_input_payload_delay_38_stateElement;
    io_input_payload_delay_40_isFull <= io_input_payload_delay_39_isFull;
    io_input_payload_delay_40_fullRound <= io_input_payload_delay_39_fullRound;
    io_input_payload_delay_40_partialRound <= io_input_payload_delay_39_partialRound;
    io_input_payload_delay_40_stateIndex <= io_input_payload_delay_39_stateIndex;
    io_input_payload_delay_40_stateSize <= io_input_payload_delay_39_stateSize;
    io_input_payload_delay_40_stateID <= io_input_payload_delay_39_stateID;
    io_input_payload_delay_40_stateElements_0 <= io_input_payload_delay_39_stateElements_0;
    io_input_payload_delay_40_stateElements_1 <= io_input_payload_delay_39_stateElements_1;
    io_input_payload_delay_40_stateElements_2 <= io_input_payload_delay_39_stateElements_2;
    io_input_payload_delay_40_stateElements_3 <= io_input_payload_delay_39_stateElements_3;
    io_input_payload_delay_40_stateElements_4 <= io_input_payload_delay_39_stateElements_4;
    io_input_payload_delay_40_stateElements_5 <= io_input_payload_delay_39_stateElements_5;
    io_input_payload_delay_40_stateElements_6 <= io_input_payload_delay_39_stateElements_6;
    io_input_payload_delay_40_stateElements_7 <= io_input_payload_delay_39_stateElements_7;
    io_input_payload_delay_40_stateElements_8 <= io_input_payload_delay_39_stateElements_8;
    io_input_payload_delay_40_stateElements_9 <= io_input_payload_delay_39_stateElements_9;
    io_input_payload_delay_40_stateElements_10 <= io_input_payload_delay_39_stateElements_10;
    io_input_payload_delay_40_stateElement <= io_input_payload_delay_39_stateElement;
    io_input_payload_delay_41_isFull <= io_input_payload_delay_40_isFull;
    io_input_payload_delay_41_fullRound <= io_input_payload_delay_40_fullRound;
    io_input_payload_delay_41_partialRound <= io_input_payload_delay_40_partialRound;
    io_input_payload_delay_41_stateIndex <= io_input_payload_delay_40_stateIndex;
    io_input_payload_delay_41_stateSize <= io_input_payload_delay_40_stateSize;
    io_input_payload_delay_41_stateID <= io_input_payload_delay_40_stateID;
    io_input_payload_delay_41_stateElements_0 <= io_input_payload_delay_40_stateElements_0;
    io_input_payload_delay_41_stateElements_1 <= io_input_payload_delay_40_stateElements_1;
    io_input_payload_delay_41_stateElements_2 <= io_input_payload_delay_40_stateElements_2;
    io_input_payload_delay_41_stateElements_3 <= io_input_payload_delay_40_stateElements_3;
    io_input_payload_delay_41_stateElements_4 <= io_input_payload_delay_40_stateElements_4;
    io_input_payload_delay_41_stateElements_5 <= io_input_payload_delay_40_stateElements_5;
    io_input_payload_delay_41_stateElements_6 <= io_input_payload_delay_40_stateElements_6;
    io_input_payload_delay_41_stateElements_7 <= io_input_payload_delay_40_stateElements_7;
    io_input_payload_delay_41_stateElements_8 <= io_input_payload_delay_40_stateElements_8;
    io_input_payload_delay_41_stateElements_9 <= io_input_payload_delay_40_stateElements_9;
    io_input_payload_delay_41_stateElements_10 <= io_input_payload_delay_40_stateElements_10;
    io_input_payload_delay_41_stateElement <= io_input_payload_delay_40_stateElement;
    io_input_payload_delay_42_isFull <= io_input_payload_delay_41_isFull;
    io_input_payload_delay_42_fullRound <= io_input_payload_delay_41_fullRound;
    io_input_payload_delay_42_partialRound <= io_input_payload_delay_41_partialRound;
    io_input_payload_delay_42_stateIndex <= io_input_payload_delay_41_stateIndex;
    io_input_payload_delay_42_stateSize <= io_input_payload_delay_41_stateSize;
    io_input_payload_delay_42_stateID <= io_input_payload_delay_41_stateID;
    io_input_payload_delay_42_stateElements_0 <= io_input_payload_delay_41_stateElements_0;
    io_input_payload_delay_42_stateElements_1 <= io_input_payload_delay_41_stateElements_1;
    io_input_payload_delay_42_stateElements_2 <= io_input_payload_delay_41_stateElements_2;
    io_input_payload_delay_42_stateElements_3 <= io_input_payload_delay_41_stateElements_3;
    io_input_payload_delay_42_stateElements_4 <= io_input_payload_delay_41_stateElements_4;
    io_input_payload_delay_42_stateElements_5 <= io_input_payload_delay_41_stateElements_5;
    io_input_payload_delay_42_stateElements_6 <= io_input_payload_delay_41_stateElements_6;
    io_input_payload_delay_42_stateElements_7 <= io_input_payload_delay_41_stateElements_7;
    io_input_payload_delay_42_stateElements_8 <= io_input_payload_delay_41_stateElements_8;
    io_input_payload_delay_42_stateElements_9 <= io_input_payload_delay_41_stateElements_9;
    io_input_payload_delay_42_stateElements_10 <= io_input_payload_delay_41_stateElements_10;
    io_input_payload_delay_42_stateElement <= io_input_payload_delay_41_stateElement;
    io_input_payload_delay_43_isFull <= io_input_payload_delay_42_isFull;
    io_input_payload_delay_43_fullRound <= io_input_payload_delay_42_fullRound;
    io_input_payload_delay_43_partialRound <= io_input_payload_delay_42_partialRound;
    io_input_payload_delay_43_stateIndex <= io_input_payload_delay_42_stateIndex;
    io_input_payload_delay_43_stateSize <= io_input_payload_delay_42_stateSize;
    io_input_payload_delay_43_stateID <= io_input_payload_delay_42_stateID;
    io_input_payload_delay_43_stateElements_0 <= io_input_payload_delay_42_stateElements_0;
    io_input_payload_delay_43_stateElements_1 <= io_input_payload_delay_42_stateElements_1;
    io_input_payload_delay_43_stateElements_2 <= io_input_payload_delay_42_stateElements_2;
    io_input_payload_delay_43_stateElements_3 <= io_input_payload_delay_42_stateElements_3;
    io_input_payload_delay_43_stateElements_4 <= io_input_payload_delay_42_stateElements_4;
    io_input_payload_delay_43_stateElements_5 <= io_input_payload_delay_42_stateElements_5;
    io_input_payload_delay_43_stateElements_6 <= io_input_payload_delay_42_stateElements_6;
    io_input_payload_delay_43_stateElements_7 <= io_input_payload_delay_42_stateElements_7;
    io_input_payload_delay_43_stateElements_8 <= io_input_payload_delay_42_stateElements_8;
    io_input_payload_delay_43_stateElements_9 <= io_input_payload_delay_42_stateElements_9;
    io_input_payload_delay_43_stateElements_10 <= io_input_payload_delay_42_stateElements_10;
    io_input_payload_delay_43_stateElement <= io_input_payload_delay_42_stateElement;
    io_input_payload_delay_44_isFull <= io_input_payload_delay_43_isFull;
    io_input_payload_delay_44_fullRound <= io_input_payload_delay_43_fullRound;
    io_input_payload_delay_44_partialRound <= io_input_payload_delay_43_partialRound;
    io_input_payload_delay_44_stateIndex <= io_input_payload_delay_43_stateIndex;
    io_input_payload_delay_44_stateSize <= io_input_payload_delay_43_stateSize;
    io_input_payload_delay_44_stateID <= io_input_payload_delay_43_stateID;
    io_input_payload_delay_44_stateElements_0 <= io_input_payload_delay_43_stateElements_0;
    io_input_payload_delay_44_stateElements_1 <= io_input_payload_delay_43_stateElements_1;
    io_input_payload_delay_44_stateElements_2 <= io_input_payload_delay_43_stateElements_2;
    io_input_payload_delay_44_stateElements_3 <= io_input_payload_delay_43_stateElements_3;
    io_input_payload_delay_44_stateElements_4 <= io_input_payload_delay_43_stateElements_4;
    io_input_payload_delay_44_stateElements_5 <= io_input_payload_delay_43_stateElements_5;
    io_input_payload_delay_44_stateElements_6 <= io_input_payload_delay_43_stateElements_6;
    io_input_payload_delay_44_stateElements_7 <= io_input_payload_delay_43_stateElements_7;
    io_input_payload_delay_44_stateElements_8 <= io_input_payload_delay_43_stateElements_8;
    io_input_payload_delay_44_stateElements_9 <= io_input_payload_delay_43_stateElements_9;
    io_input_payload_delay_44_stateElements_10 <= io_input_payload_delay_43_stateElements_10;
    io_input_payload_delay_44_stateElement <= io_input_payload_delay_43_stateElement;
    io_input_payload_delay_45_isFull <= io_input_payload_delay_44_isFull;
    io_input_payload_delay_45_fullRound <= io_input_payload_delay_44_fullRound;
    io_input_payload_delay_45_partialRound <= io_input_payload_delay_44_partialRound;
    io_input_payload_delay_45_stateIndex <= io_input_payload_delay_44_stateIndex;
    io_input_payload_delay_45_stateSize <= io_input_payload_delay_44_stateSize;
    io_input_payload_delay_45_stateID <= io_input_payload_delay_44_stateID;
    io_input_payload_delay_45_stateElements_0 <= io_input_payload_delay_44_stateElements_0;
    io_input_payload_delay_45_stateElements_1 <= io_input_payload_delay_44_stateElements_1;
    io_input_payload_delay_45_stateElements_2 <= io_input_payload_delay_44_stateElements_2;
    io_input_payload_delay_45_stateElements_3 <= io_input_payload_delay_44_stateElements_3;
    io_input_payload_delay_45_stateElements_4 <= io_input_payload_delay_44_stateElements_4;
    io_input_payload_delay_45_stateElements_5 <= io_input_payload_delay_44_stateElements_5;
    io_input_payload_delay_45_stateElements_6 <= io_input_payload_delay_44_stateElements_6;
    io_input_payload_delay_45_stateElements_7 <= io_input_payload_delay_44_stateElements_7;
    io_input_payload_delay_45_stateElements_8 <= io_input_payload_delay_44_stateElements_8;
    io_input_payload_delay_45_stateElements_9 <= io_input_payload_delay_44_stateElements_9;
    io_input_payload_delay_45_stateElements_10 <= io_input_payload_delay_44_stateElements_10;
    io_input_payload_delay_45_stateElement <= io_input_payload_delay_44_stateElement;
    io_input_payload_delay_46_isFull <= io_input_payload_delay_45_isFull;
    io_input_payload_delay_46_fullRound <= io_input_payload_delay_45_fullRound;
    io_input_payload_delay_46_partialRound <= io_input_payload_delay_45_partialRound;
    io_input_payload_delay_46_stateIndex <= io_input_payload_delay_45_stateIndex;
    io_input_payload_delay_46_stateSize <= io_input_payload_delay_45_stateSize;
    io_input_payload_delay_46_stateID <= io_input_payload_delay_45_stateID;
    io_input_payload_delay_46_stateElements_0 <= io_input_payload_delay_45_stateElements_0;
    io_input_payload_delay_46_stateElements_1 <= io_input_payload_delay_45_stateElements_1;
    io_input_payload_delay_46_stateElements_2 <= io_input_payload_delay_45_stateElements_2;
    io_input_payload_delay_46_stateElements_3 <= io_input_payload_delay_45_stateElements_3;
    io_input_payload_delay_46_stateElements_4 <= io_input_payload_delay_45_stateElements_4;
    io_input_payload_delay_46_stateElements_5 <= io_input_payload_delay_45_stateElements_5;
    io_input_payload_delay_46_stateElements_6 <= io_input_payload_delay_45_stateElements_6;
    io_input_payload_delay_46_stateElements_7 <= io_input_payload_delay_45_stateElements_7;
    io_input_payload_delay_46_stateElements_8 <= io_input_payload_delay_45_stateElements_8;
    io_input_payload_delay_46_stateElements_9 <= io_input_payload_delay_45_stateElements_9;
    io_input_payload_delay_46_stateElements_10 <= io_input_payload_delay_45_stateElements_10;
    io_input_payload_delay_46_stateElement <= io_input_payload_delay_45_stateElement;
    io_input_payload_delay_47_isFull <= io_input_payload_delay_46_isFull;
    io_input_payload_delay_47_fullRound <= io_input_payload_delay_46_fullRound;
    io_input_payload_delay_47_partialRound <= io_input_payload_delay_46_partialRound;
    io_input_payload_delay_47_stateIndex <= io_input_payload_delay_46_stateIndex;
    io_input_payload_delay_47_stateSize <= io_input_payload_delay_46_stateSize;
    io_input_payload_delay_47_stateID <= io_input_payload_delay_46_stateID;
    io_input_payload_delay_47_stateElements_0 <= io_input_payload_delay_46_stateElements_0;
    io_input_payload_delay_47_stateElements_1 <= io_input_payload_delay_46_stateElements_1;
    io_input_payload_delay_47_stateElements_2 <= io_input_payload_delay_46_stateElements_2;
    io_input_payload_delay_47_stateElements_3 <= io_input_payload_delay_46_stateElements_3;
    io_input_payload_delay_47_stateElements_4 <= io_input_payload_delay_46_stateElements_4;
    io_input_payload_delay_47_stateElements_5 <= io_input_payload_delay_46_stateElements_5;
    io_input_payload_delay_47_stateElements_6 <= io_input_payload_delay_46_stateElements_6;
    io_input_payload_delay_47_stateElements_7 <= io_input_payload_delay_46_stateElements_7;
    io_input_payload_delay_47_stateElements_8 <= io_input_payload_delay_46_stateElements_8;
    io_input_payload_delay_47_stateElements_9 <= io_input_payload_delay_46_stateElements_9;
    io_input_payload_delay_47_stateElements_10 <= io_input_payload_delay_46_stateElements_10;
    io_input_payload_delay_47_stateElement <= io_input_payload_delay_46_stateElement;
    io_input_payload_delay_48_isFull <= io_input_payload_delay_47_isFull;
    io_input_payload_delay_48_fullRound <= io_input_payload_delay_47_fullRound;
    io_input_payload_delay_48_partialRound <= io_input_payload_delay_47_partialRound;
    io_input_payload_delay_48_stateIndex <= io_input_payload_delay_47_stateIndex;
    io_input_payload_delay_48_stateSize <= io_input_payload_delay_47_stateSize;
    io_input_payload_delay_48_stateID <= io_input_payload_delay_47_stateID;
    io_input_payload_delay_48_stateElements_0 <= io_input_payload_delay_47_stateElements_0;
    io_input_payload_delay_48_stateElements_1 <= io_input_payload_delay_47_stateElements_1;
    io_input_payload_delay_48_stateElements_2 <= io_input_payload_delay_47_stateElements_2;
    io_input_payload_delay_48_stateElements_3 <= io_input_payload_delay_47_stateElements_3;
    io_input_payload_delay_48_stateElements_4 <= io_input_payload_delay_47_stateElements_4;
    io_input_payload_delay_48_stateElements_5 <= io_input_payload_delay_47_stateElements_5;
    io_input_payload_delay_48_stateElements_6 <= io_input_payload_delay_47_stateElements_6;
    io_input_payload_delay_48_stateElements_7 <= io_input_payload_delay_47_stateElements_7;
    io_input_payload_delay_48_stateElements_8 <= io_input_payload_delay_47_stateElements_8;
    io_input_payload_delay_48_stateElements_9 <= io_input_payload_delay_47_stateElements_9;
    io_input_payload_delay_48_stateElements_10 <= io_input_payload_delay_47_stateElements_10;
    io_input_payload_delay_48_stateElement <= io_input_payload_delay_47_stateElement;
    io_input_payload_delay_49_isFull <= io_input_payload_delay_48_isFull;
    io_input_payload_delay_49_fullRound <= io_input_payload_delay_48_fullRound;
    io_input_payload_delay_49_partialRound <= io_input_payload_delay_48_partialRound;
    io_input_payload_delay_49_stateIndex <= io_input_payload_delay_48_stateIndex;
    io_input_payload_delay_49_stateSize <= io_input_payload_delay_48_stateSize;
    io_input_payload_delay_49_stateID <= io_input_payload_delay_48_stateID;
    io_input_payload_delay_49_stateElements_0 <= io_input_payload_delay_48_stateElements_0;
    io_input_payload_delay_49_stateElements_1 <= io_input_payload_delay_48_stateElements_1;
    io_input_payload_delay_49_stateElements_2 <= io_input_payload_delay_48_stateElements_2;
    io_input_payload_delay_49_stateElements_3 <= io_input_payload_delay_48_stateElements_3;
    io_input_payload_delay_49_stateElements_4 <= io_input_payload_delay_48_stateElements_4;
    io_input_payload_delay_49_stateElements_5 <= io_input_payload_delay_48_stateElements_5;
    io_input_payload_delay_49_stateElements_6 <= io_input_payload_delay_48_stateElements_6;
    io_input_payload_delay_49_stateElements_7 <= io_input_payload_delay_48_stateElements_7;
    io_input_payload_delay_49_stateElements_8 <= io_input_payload_delay_48_stateElements_8;
    io_input_payload_delay_49_stateElements_9 <= io_input_payload_delay_48_stateElements_9;
    io_input_payload_delay_49_stateElements_10 <= io_input_payload_delay_48_stateElements_10;
    io_input_payload_delay_49_stateElement <= io_input_payload_delay_48_stateElement;
    io_input_payload_delay_50_isFull <= io_input_payload_delay_49_isFull;
    io_input_payload_delay_50_fullRound <= io_input_payload_delay_49_fullRound;
    io_input_payload_delay_50_partialRound <= io_input_payload_delay_49_partialRound;
    io_input_payload_delay_50_stateIndex <= io_input_payload_delay_49_stateIndex;
    io_input_payload_delay_50_stateSize <= io_input_payload_delay_49_stateSize;
    io_input_payload_delay_50_stateID <= io_input_payload_delay_49_stateID;
    io_input_payload_delay_50_stateElements_0 <= io_input_payload_delay_49_stateElements_0;
    io_input_payload_delay_50_stateElements_1 <= io_input_payload_delay_49_stateElements_1;
    io_input_payload_delay_50_stateElements_2 <= io_input_payload_delay_49_stateElements_2;
    io_input_payload_delay_50_stateElements_3 <= io_input_payload_delay_49_stateElements_3;
    io_input_payload_delay_50_stateElements_4 <= io_input_payload_delay_49_stateElements_4;
    io_input_payload_delay_50_stateElements_5 <= io_input_payload_delay_49_stateElements_5;
    io_input_payload_delay_50_stateElements_6 <= io_input_payload_delay_49_stateElements_6;
    io_input_payload_delay_50_stateElements_7 <= io_input_payload_delay_49_stateElements_7;
    io_input_payload_delay_50_stateElements_8 <= io_input_payload_delay_49_stateElements_8;
    io_input_payload_delay_50_stateElements_9 <= io_input_payload_delay_49_stateElements_9;
    io_input_payload_delay_50_stateElements_10 <= io_input_payload_delay_49_stateElements_10;
    io_input_payload_delay_50_stateElement <= io_input_payload_delay_49_stateElement;
    io_input_payload_delay_51_isFull <= io_input_payload_delay_50_isFull;
    io_input_payload_delay_51_fullRound <= io_input_payload_delay_50_fullRound;
    io_input_payload_delay_51_partialRound <= io_input_payload_delay_50_partialRound;
    io_input_payload_delay_51_stateIndex <= io_input_payload_delay_50_stateIndex;
    io_input_payload_delay_51_stateSize <= io_input_payload_delay_50_stateSize;
    io_input_payload_delay_51_stateID <= io_input_payload_delay_50_stateID;
    io_input_payload_delay_51_stateElements_0 <= io_input_payload_delay_50_stateElements_0;
    io_input_payload_delay_51_stateElements_1 <= io_input_payload_delay_50_stateElements_1;
    io_input_payload_delay_51_stateElements_2 <= io_input_payload_delay_50_stateElements_2;
    io_input_payload_delay_51_stateElements_3 <= io_input_payload_delay_50_stateElements_3;
    io_input_payload_delay_51_stateElements_4 <= io_input_payload_delay_50_stateElements_4;
    io_input_payload_delay_51_stateElements_5 <= io_input_payload_delay_50_stateElements_5;
    io_input_payload_delay_51_stateElements_6 <= io_input_payload_delay_50_stateElements_6;
    io_input_payload_delay_51_stateElements_7 <= io_input_payload_delay_50_stateElements_7;
    io_input_payload_delay_51_stateElements_8 <= io_input_payload_delay_50_stateElements_8;
    io_input_payload_delay_51_stateElements_9 <= io_input_payload_delay_50_stateElements_9;
    io_input_payload_delay_51_stateElements_10 <= io_input_payload_delay_50_stateElements_10;
    io_input_payload_delay_51_stateElement <= io_input_payload_delay_50_stateElement;
    io_input_payload_delay_52_isFull <= io_input_payload_delay_51_isFull;
    io_input_payload_delay_52_fullRound <= io_input_payload_delay_51_fullRound;
    io_input_payload_delay_52_partialRound <= io_input_payload_delay_51_partialRound;
    io_input_payload_delay_52_stateIndex <= io_input_payload_delay_51_stateIndex;
    io_input_payload_delay_52_stateSize <= io_input_payload_delay_51_stateSize;
    io_input_payload_delay_52_stateID <= io_input_payload_delay_51_stateID;
    io_input_payload_delay_52_stateElements_0 <= io_input_payload_delay_51_stateElements_0;
    io_input_payload_delay_52_stateElements_1 <= io_input_payload_delay_51_stateElements_1;
    io_input_payload_delay_52_stateElements_2 <= io_input_payload_delay_51_stateElements_2;
    io_input_payload_delay_52_stateElements_3 <= io_input_payload_delay_51_stateElements_3;
    io_input_payload_delay_52_stateElements_4 <= io_input_payload_delay_51_stateElements_4;
    io_input_payload_delay_52_stateElements_5 <= io_input_payload_delay_51_stateElements_5;
    io_input_payload_delay_52_stateElements_6 <= io_input_payload_delay_51_stateElements_6;
    io_input_payload_delay_52_stateElements_7 <= io_input_payload_delay_51_stateElements_7;
    io_input_payload_delay_52_stateElements_8 <= io_input_payload_delay_51_stateElements_8;
    io_input_payload_delay_52_stateElements_9 <= io_input_payload_delay_51_stateElements_9;
    io_input_payload_delay_52_stateElements_10 <= io_input_payload_delay_51_stateElements_10;
    io_input_payload_delay_52_stateElement <= io_input_payload_delay_51_stateElement;
    io_input_payload_delay_53_isFull <= io_input_payload_delay_52_isFull;
    io_input_payload_delay_53_fullRound <= io_input_payload_delay_52_fullRound;
    io_input_payload_delay_53_partialRound <= io_input_payload_delay_52_partialRound;
    io_input_payload_delay_53_stateIndex <= io_input_payload_delay_52_stateIndex;
    io_input_payload_delay_53_stateSize <= io_input_payload_delay_52_stateSize;
    io_input_payload_delay_53_stateID <= io_input_payload_delay_52_stateID;
    io_input_payload_delay_53_stateElements_0 <= io_input_payload_delay_52_stateElements_0;
    io_input_payload_delay_53_stateElements_1 <= io_input_payload_delay_52_stateElements_1;
    io_input_payload_delay_53_stateElements_2 <= io_input_payload_delay_52_stateElements_2;
    io_input_payload_delay_53_stateElements_3 <= io_input_payload_delay_52_stateElements_3;
    io_input_payload_delay_53_stateElements_4 <= io_input_payload_delay_52_stateElements_4;
    io_input_payload_delay_53_stateElements_5 <= io_input_payload_delay_52_stateElements_5;
    io_input_payload_delay_53_stateElements_6 <= io_input_payload_delay_52_stateElements_6;
    io_input_payload_delay_53_stateElements_7 <= io_input_payload_delay_52_stateElements_7;
    io_input_payload_delay_53_stateElements_8 <= io_input_payload_delay_52_stateElements_8;
    io_input_payload_delay_53_stateElements_9 <= io_input_payload_delay_52_stateElements_9;
    io_input_payload_delay_53_stateElements_10 <= io_input_payload_delay_52_stateElements_10;
    io_input_payload_delay_53_stateElement <= io_input_payload_delay_52_stateElement;
    io_input_payload_delay_54_isFull <= io_input_payload_delay_53_isFull;
    io_input_payload_delay_54_fullRound <= io_input_payload_delay_53_fullRound;
    io_input_payload_delay_54_partialRound <= io_input_payload_delay_53_partialRound;
    io_input_payload_delay_54_stateIndex <= io_input_payload_delay_53_stateIndex;
    io_input_payload_delay_54_stateSize <= io_input_payload_delay_53_stateSize;
    io_input_payload_delay_54_stateID <= io_input_payload_delay_53_stateID;
    io_input_payload_delay_54_stateElements_0 <= io_input_payload_delay_53_stateElements_0;
    io_input_payload_delay_54_stateElements_1 <= io_input_payload_delay_53_stateElements_1;
    io_input_payload_delay_54_stateElements_2 <= io_input_payload_delay_53_stateElements_2;
    io_input_payload_delay_54_stateElements_3 <= io_input_payload_delay_53_stateElements_3;
    io_input_payload_delay_54_stateElements_4 <= io_input_payload_delay_53_stateElements_4;
    io_input_payload_delay_54_stateElements_5 <= io_input_payload_delay_53_stateElements_5;
    io_input_payload_delay_54_stateElements_6 <= io_input_payload_delay_53_stateElements_6;
    io_input_payload_delay_54_stateElements_7 <= io_input_payload_delay_53_stateElements_7;
    io_input_payload_delay_54_stateElements_8 <= io_input_payload_delay_53_stateElements_8;
    io_input_payload_delay_54_stateElements_9 <= io_input_payload_delay_53_stateElements_9;
    io_input_payload_delay_54_stateElements_10 <= io_input_payload_delay_53_stateElements_10;
    io_input_payload_delay_54_stateElement <= io_input_payload_delay_53_stateElement;
    io_input_payload_delay_55_isFull <= io_input_payload_delay_54_isFull;
    io_input_payload_delay_55_fullRound <= io_input_payload_delay_54_fullRound;
    io_input_payload_delay_55_partialRound <= io_input_payload_delay_54_partialRound;
    io_input_payload_delay_55_stateIndex <= io_input_payload_delay_54_stateIndex;
    io_input_payload_delay_55_stateSize <= io_input_payload_delay_54_stateSize;
    io_input_payload_delay_55_stateID <= io_input_payload_delay_54_stateID;
    io_input_payload_delay_55_stateElements_0 <= io_input_payload_delay_54_stateElements_0;
    io_input_payload_delay_55_stateElements_1 <= io_input_payload_delay_54_stateElements_1;
    io_input_payload_delay_55_stateElements_2 <= io_input_payload_delay_54_stateElements_2;
    io_input_payload_delay_55_stateElements_3 <= io_input_payload_delay_54_stateElements_3;
    io_input_payload_delay_55_stateElements_4 <= io_input_payload_delay_54_stateElements_4;
    io_input_payload_delay_55_stateElements_5 <= io_input_payload_delay_54_stateElements_5;
    io_input_payload_delay_55_stateElements_6 <= io_input_payload_delay_54_stateElements_6;
    io_input_payload_delay_55_stateElements_7 <= io_input_payload_delay_54_stateElements_7;
    io_input_payload_delay_55_stateElements_8 <= io_input_payload_delay_54_stateElements_8;
    io_input_payload_delay_55_stateElements_9 <= io_input_payload_delay_54_stateElements_9;
    io_input_payload_delay_55_stateElements_10 <= io_input_payload_delay_54_stateElements_10;
    io_input_payload_delay_55_stateElement <= io_input_payload_delay_54_stateElement;
    io_input_payload_delay_56_isFull <= io_input_payload_delay_55_isFull;
    io_input_payload_delay_56_fullRound <= io_input_payload_delay_55_fullRound;
    io_input_payload_delay_56_partialRound <= io_input_payload_delay_55_partialRound;
    io_input_payload_delay_56_stateIndex <= io_input_payload_delay_55_stateIndex;
    io_input_payload_delay_56_stateSize <= io_input_payload_delay_55_stateSize;
    io_input_payload_delay_56_stateID <= io_input_payload_delay_55_stateID;
    io_input_payload_delay_56_stateElements_0 <= io_input_payload_delay_55_stateElements_0;
    io_input_payload_delay_56_stateElements_1 <= io_input_payload_delay_55_stateElements_1;
    io_input_payload_delay_56_stateElements_2 <= io_input_payload_delay_55_stateElements_2;
    io_input_payload_delay_56_stateElements_3 <= io_input_payload_delay_55_stateElements_3;
    io_input_payload_delay_56_stateElements_4 <= io_input_payload_delay_55_stateElements_4;
    io_input_payload_delay_56_stateElements_5 <= io_input_payload_delay_55_stateElements_5;
    io_input_payload_delay_56_stateElements_6 <= io_input_payload_delay_55_stateElements_6;
    io_input_payload_delay_56_stateElements_7 <= io_input_payload_delay_55_stateElements_7;
    io_input_payload_delay_56_stateElements_8 <= io_input_payload_delay_55_stateElements_8;
    io_input_payload_delay_56_stateElements_9 <= io_input_payload_delay_55_stateElements_9;
    io_input_payload_delay_56_stateElements_10 <= io_input_payload_delay_55_stateElements_10;
    io_input_payload_delay_56_stateElement <= io_input_payload_delay_55_stateElement;
    io_input_payload_delay_57_isFull <= io_input_payload_delay_56_isFull;
    io_input_payload_delay_57_fullRound <= io_input_payload_delay_56_fullRound;
    io_input_payload_delay_57_partialRound <= io_input_payload_delay_56_partialRound;
    io_input_payload_delay_57_stateIndex <= io_input_payload_delay_56_stateIndex;
    io_input_payload_delay_57_stateSize <= io_input_payload_delay_56_stateSize;
    io_input_payload_delay_57_stateID <= io_input_payload_delay_56_stateID;
    io_input_payload_delay_57_stateElements_0 <= io_input_payload_delay_56_stateElements_0;
    io_input_payload_delay_57_stateElements_1 <= io_input_payload_delay_56_stateElements_1;
    io_input_payload_delay_57_stateElements_2 <= io_input_payload_delay_56_stateElements_2;
    io_input_payload_delay_57_stateElements_3 <= io_input_payload_delay_56_stateElements_3;
    io_input_payload_delay_57_stateElements_4 <= io_input_payload_delay_56_stateElements_4;
    io_input_payload_delay_57_stateElements_5 <= io_input_payload_delay_56_stateElements_5;
    io_input_payload_delay_57_stateElements_6 <= io_input_payload_delay_56_stateElements_6;
    io_input_payload_delay_57_stateElements_7 <= io_input_payload_delay_56_stateElements_7;
    io_input_payload_delay_57_stateElements_8 <= io_input_payload_delay_56_stateElements_8;
    io_input_payload_delay_57_stateElements_9 <= io_input_payload_delay_56_stateElements_9;
    io_input_payload_delay_57_stateElements_10 <= io_input_payload_delay_56_stateElements_10;
    io_input_payload_delay_57_stateElement <= io_input_payload_delay_56_stateElement;
    io_input_payload_delay_58_isFull <= io_input_payload_delay_57_isFull;
    io_input_payload_delay_58_fullRound <= io_input_payload_delay_57_fullRound;
    io_input_payload_delay_58_partialRound <= io_input_payload_delay_57_partialRound;
    io_input_payload_delay_58_stateIndex <= io_input_payload_delay_57_stateIndex;
    io_input_payload_delay_58_stateSize <= io_input_payload_delay_57_stateSize;
    io_input_payload_delay_58_stateID <= io_input_payload_delay_57_stateID;
    io_input_payload_delay_58_stateElements_0 <= io_input_payload_delay_57_stateElements_0;
    io_input_payload_delay_58_stateElements_1 <= io_input_payload_delay_57_stateElements_1;
    io_input_payload_delay_58_stateElements_2 <= io_input_payload_delay_57_stateElements_2;
    io_input_payload_delay_58_stateElements_3 <= io_input_payload_delay_57_stateElements_3;
    io_input_payload_delay_58_stateElements_4 <= io_input_payload_delay_57_stateElements_4;
    io_input_payload_delay_58_stateElements_5 <= io_input_payload_delay_57_stateElements_5;
    io_input_payload_delay_58_stateElements_6 <= io_input_payload_delay_57_stateElements_6;
    io_input_payload_delay_58_stateElements_7 <= io_input_payload_delay_57_stateElements_7;
    io_input_payload_delay_58_stateElements_8 <= io_input_payload_delay_57_stateElements_8;
    io_input_payload_delay_58_stateElements_9 <= io_input_payload_delay_57_stateElements_9;
    io_input_payload_delay_58_stateElements_10 <= io_input_payload_delay_57_stateElements_10;
    io_input_payload_delay_58_stateElement <= io_input_payload_delay_57_stateElement;
    io_input_payload_delay_59_isFull <= io_input_payload_delay_58_isFull;
    io_input_payload_delay_59_fullRound <= io_input_payload_delay_58_fullRound;
    io_input_payload_delay_59_partialRound <= io_input_payload_delay_58_partialRound;
    io_input_payload_delay_59_stateIndex <= io_input_payload_delay_58_stateIndex;
    io_input_payload_delay_59_stateSize <= io_input_payload_delay_58_stateSize;
    io_input_payload_delay_59_stateID <= io_input_payload_delay_58_stateID;
    io_input_payload_delay_59_stateElements_0 <= io_input_payload_delay_58_stateElements_0;
    io_input_payload_delay_59_stateElements_1 <= io_input_payload_delay_58_stateElements_1;
    io_input_payload_delay_59_stateElements_2 <= io_input_payload_delay_58_stateElements_2;
    io_input_payload_delay_59_stateElements_3 <= io_input_payload_delay_58_stateElements_3;
    io_input_payload_delay_59_stateElements_4 <= io_input_payload_delay_58_stateElements_4;
    io_input_payload_delay_59_stateElements_5 <= io_input_payload_delay_58_stateElements_5;
    io_input_payload_delay_59_stateElements_6 <= io_input_payload_delay_58_stateElements_6;
    io_input_payload_delay_59_stateElements_7 <= io_input_payload_delay_58_stateElements_7;
    io_input_payload_delay_59_stateElements_8 <= io_input_payload_delay_58_stateElements_8;
    io_input_payload_delay_59_stateElements_9 <= io_input_payload_delay_58_stateElements_9;
    io_input_payload_delay_59_stateElements_10 <= io_input_payload_delay_58_stateElements_10;
    io_input_payload_delay_59_stateElement <= io_input_payload_delay_58_stateElement;
    io_input_payload_delay_60_isFull <= io_input_payload_delay_59_isFull;
    io_input_payload_delay_60_fullRound <= io_input_payload_delay_59_fullRound;
    io_input_payload_delay_60_partialRound <= io_input_payload_delay_59_partialRound;
    io_input_payload_delay_60_stateIndex <= io_input_payload_delay_59_stateIndex;
    io_input_payload_delay_60_stateSize <= io_input_payload_delay_59_stateSize;
    io_input_payload_delay_60_stateID <= io_input_payload_delay_59_stateID;
    io_input_payload_delay_60_stateElements_0 <= io_input_payload_delay_59_stateElements_0;
    io_input_payload_delay_60_stateElements_1 <= io_input_payload_delay_59_stateElements_1;
    io_input_payload_delay_60_stateElements_2 <= io_input_payload_delay_59_stateElements_2;
    io_input_payload_delay_60_stateElements_3 <= io_input_payload_delay_59_stateElements_3;
    io_input_payload_delay_60_stateElements_4 <= io_input_payload_delay_59_stateElements_4;
    io_input_payload_delay_60_stateElements_5 <= io_input_payload_delay_59_stateElements_5;
    io_input_payload_delay_60_stateElements_6 <= io_input_payload_delay_59_stateElements_6;
    io_input_payload_delay_60_stateElements_7 <= io_input_payload_delay_59_stateElements_7;
    io_input_payload_delay_60_stateElements_8 <= io_input_payload_delay_59_stateElements_8;
    io_input_payload_delay_60_stateElements_9 <= io_input_payload_delay_59_stateElements_9;
    io_input_payload_delay_60_stateElements_10 <= io_input_payload_delay_59_stateElements_10;
    io_input_payload_delay_60_stateElement <= io_input_payload_delay_59_stateElement;
    io_input_payload_delay_61_isFull <= io_input_payload_delay_60_isFull;
    io_input_payload_delay_61_fullRound <= io_input_payload_delay_60_fullRound;
    io_input_payload_delay_61_partialRound <= io_input_payload_delay_60_partialRound;
    io_input_payload_delay_61_stateIndex <= io_input_payload_delay_60_stateIndex;
    io_input_payload_delay_61_stateSize <= io_input_payload_delay_60_stateSize;
    io_input_payload_delay_61_stateID <= io_input_payload_delay_60_stateID;
    io_input_payload_delay_61_stateElements_0 <= io_input_payload_delay_60_stateElements_0;
    io_input_payload_delay_61_stateElements_1 <= io_input_payload_delay_60_stateElements_1;
    io_input_payload_delay_61_stateElements_2 <= io_input_payload_delay_60_stateElements_2;
    io_input_payload_delay_61_stateElements_3 <= io_input_payload_delay_60_stateElements_3;
    io_input_payload_delay_61_stateElements_4 <= io_input_payload_delay_60_stateElements_4;
    io_input_payload_delay_61_stateElements_5 <= io_input_payload_delay_60_stateElements_5;
    io_input_payload_delay_61_stateElements_6 <= io_input_payload_delay_60_stateElements_6;
    io_input_payload_delay_61_stateElements_7 <= io_input_payload_delay_60_stateElements_7;
    io_input_payload_delay_61_stateElements_8 <= io_input_payload_delay_60_stateElements_8;
    io_input_payload_delay_61_stateElements_9 <= io_input_payload_delay_60_stateElements_9;
    io_input_payload_delay_61_stateElements_10 <= io_input_payload_delay_60_stateElements_10;
    io_input_payload_delay_61_stateElement <= io_input_payload_delay_60_stateElement;
    io_input_payload_delay_62_isFull <= io_input_payload_delay_61_isFull;
    io_input_payload_delay_62_fullRound <= io_input_payload_delay_61_fullRound;
    io_input_payload_delay_62_partialRound <= io_input_payload_delay_61_partialRound;
    io_input_payload_delay_62_stateIndex <= io_input_payload_delay_61_stateIndex;
    io_input_payload_delay_62_stateSize <= io_input_payload_delay_61_stateSize;
    io_input_payload_delay_62_stateID <= io_input_payload_delay_61_stateID;
    io_input_payload_delay_62_stateElements_0 <= io_input_payload_delay_61_stateElements_0;
    io_input_payload_delay_62_stateElements_1 <= io_input_payload_delay_61_stateElements_1;
    io_input_payload_delay_62_stateElements_2 <= io_input_payload_delay_61_stateElements_2;
    io_input_payload_delay_62_stateElements_3 <= io_input_payload_delay_61_stateElements_3;
    io_input_payload_delay_62_stateElements_4 <= io_input_payload_delay_61_stateElements_4;
    io_input_payload_delay_62_stateElements_5 <= io_input_payload_delay_61_stateElements_5;
    io_input_payload_delay_62_stateElements_6 <= io_input_payload_delay_61_stateElements_6;
    io_input_payload_delay_62_stateElements_7 <= io_input_payload_delay_61_stateElements_7;
    io_input_payload_delay_62_stateElements_8 <= io_input_payload_delay_61_stateElements_8;
    io_input_payload_delay_62_stateElements_9 <= io_input_payload_delay_61_stateElements_9;
    io_input_payload_delay_62_stateElements_10 <= io_input_payload_delay_61_stateElements_10;
    io_input_payload_delay_62_stateElement <= io_input_payload_delay_61_stateElement;
    io_input_payload_delay_63_isFull <= io_input_payload_delay_62_isFull;
    io_input_payload_delay_63_fullRound <= io_input_payload_delay_62_fullRound;
    io_input_payload_delay_63_partialRound <= io_input_payload_delay_62_partialRound;
    io_input_payload_delay_63_stateIndex <= io_input_payload_delay_62_stateIndex;
    io_input_payload_delay_63_stateSize <= io_input_payload_delay_62_stateSize;
    io_input_payload_delay_63_stateID <= io_input_payload_delay_62_stateID;
    io_input_payload_delay_63_stateElements_0 <= io_input_payload_delay_62_stateElements_0;
    io_input_payload_delay_63_stateElements_1 <= io_input_payload_delay_62_stateElements_1;
    io_input_payload_delay_63_stateElements_2 <= io_input_payload_delay_62_stateElements_2;
    io_input_payload_delay_63_stateElements_3 <= io_input_payload_delay_62_stateElements_3;
    io_input_payload_delay_63_stateElements_4 <= io_input_payload_delay_62_stateElements_4;
    io_input_payload_delay_63_stateElements_5 <= io_input_payload_delay_62_stateElements_5;
    io_input_payload_delay_63_stateElements_6 <= io_input_payload_delay_62_stateElements_6;
    io_input_payload_delay_63_stateElements_7 <= io_input_payload_delay_62_stateElements_7;
    io_input_payload_delay_63_stateElements_8 <= io_input_payload_delay_62_stateElements_8;
    io_input_payload_delay_63_stateElements_9 <= io_input_payload_delay_62_stateElements_9;
    io_input_payload_delay_63_stateElements_10 <= io_input_payload_delay_62_stateElements_10;
    io_input_payload_delay_63_stateElement <= io_input_payload_delay_62_stateElement;
    io_input_payload_delay_64_isFull <= io_input_payload_delay_63_isFull;
    io_input_payload_delay_64_fullRound <= io_input_payload_delay_63_fullRound;
    io_input_payload_delay_64_partialRound <= io_input_payload_delay_63_partialRound;
    io_input_payload_delay_64_stateIndex <= io_input_payload_delay_63_stateIndex;
    io_input_payload_delay_64_stateSize <= io_input_payload_delay_63_stateSize;
    io_input_payload_delay_64_stateID <= io_input_payload_delay_63_stateID;
    io_input_payload_delay_64_stateElements_0 <= io_input_payload_delay_63_stateElements_0;
    io_input_payload_delay_64_stateElements_1 <= io_input_payload_delay_63_stateElements_1;
    io_input_payload_delay_64_stateElements_2 <= io_input_payload_delay_63_stateElements_2;
    io_input_payload_delay_64_stateElements_3 <= io_input_payload_delay_63_stateElements_3;
    io_input_payload_delay_64_stateElements_4 <= io_input_payload_delay_63_stateElements_4;
    io_input_payload_delay_64_stateElements_5 <= io_input_payload_delay_63_stateElements_5;
    io_input_payload_delay_64_stateElements_6 <= io_input_payload_delay_63_stateElements_6;
    io_input_payload_delay_64_stateElements_7 <= io_input_payload_delay_63_stateElements_7;
    io_input_payload_delay_64_stateElements_8 <= io_input_payload_delay_63_stateElements_8;
    io_input_payload_delay_64_stateElements_9 <= io_input_payload_delay_63_stateElements_9;
    io_input_payload_delay_64_stateElements_10 <= io_input_payload_delay_63_stateElements_10;
    io_input_payload_delay_64_stateElement <= io_input_payload_delay_63_stateElement;
    io_input_payload_delay_65_isFull <= io_input_payload_delay_64_isFull;
    io_input_payload_delay_65_fullRound <= io_input_payload_delay_64_fullRound;
    io_input_payload_delay_65_partialRound <= io_input_payload_delay_64_partialRound;
    io_input_payload_delay_65_stateIndex <= io_input_payload_delay_64_stateIndex;
    io_input_payload_delay_65_stateSize <= io_input_payload_delay_64_stateSize;
    io_input_payload_delay_65_stateID <= io_input_payload_delay_64_stateID;
    io_input_payload_delay_65_stateElements_0 <= io_input_payload_delay_64_stateElements_0;
    io_input_payload_delay_65_stateElements_1 <= io_input_payload_delay_64_stateElements_1;
    io_input_payload_delay_65_stateElements_2 <= io_input_payload_delay_64_stateElements_2;
    io_input_payload_delay_65_stateElements_3 <= io_input_payload_delay_64_stateElements_3;
    io_input_payload_delay_65_stateElements_4 <= io_input_payload_delay_64_stateElements_4;
    io_input_payload_delay_65_stateElements_5 <= io_input_payload_delay_64_stateElements_5;
    io_input_payload_delay_65_stateElements_6 <= io_input_payload_delay_64_stateElements_6;
    io_input_payload_delay_65_stateElements_7 <= io_input_payload_delay_64_stateElements_7;
    io_input_payload_delay_65_stateElements_8 <= io_input_payload_delay_64_stateElements_8;
    io_input_payload_delay_65_stateElements_9 <= io_input_payload_delay_64_stateElements_9;
    io_input_payload_delay_65_stateElements_10 <= io_input_payload_delay_64_stateElements_10;
    io_input_payload_delay_65_stateElement <= io_input_payload_delay_64_stateElement;
    io_input_payload_delay_66_isFull <= io_input_payload_delay_65_isFull;
    io_input_payload_delay_66_fullRound <= io_input_payload_delay_65_fullRound;
    io_input_payload_delay_66_partialRound <= io_input_payload_delay_65_partialRound;
    io_input_payload_delay_66_stateIndex <= io_input_payload_delay_65_stateIndex;
    io_input_payload_delay_66_stateSize <= io_input_payload_delay_65_stateSize;
    io_input_payload_delay_66_stateID <= io_input_payload_delay_65_stateID;
    io_input_payload_delay_66_stateElements_0 <= io_input_payload_delay_65_stateElements_0;
    io_input_payload_delay_66_stateElements_1 <= io_input_payload_delay_65_stateElements_1;
    io_input_payload_delay_66_stateElements_2 <= io_input_payload_delay_65_stateElements_2;
    io_input_payload_delay_66_stateElements_3 <= io_input_payload_delay_65_stateElements_3;
    io_input_payload_delay_66_stateElements_4 <= io_input_payload_delay_65_stateElements_4;
    io_input_payload_delay_66_stateElements_5 <= io_input_payload_delay_65_stateElements_5;
    io_input_payload_delay_66_stateElements_6 <= io_input_payload_delay_65_stateElements_6;
    io_input_payload_delay_66_stateElements_7 <= io_input_payload_delay_65_stateElements_7;
    io_input_payload_delay_66_stateElements_8 <= io_input_payload_delay_65_stateElements_8;
    io_input_payload_delay_66_stateElements_9 <= io_input_payload_delay_65_stateElements_9;
    io_input_payload_delay_66_stateElements_10 <= io_input_payload_delay_65_stateElements_10;
    io_input_payload_delay_66_stateElement <= io_input_payload_delay_65_stateElement;
    io_input_payload_delay_67_isFull <= io_input_payload_delay_66_isFull;
    io_input_payload_delay_67_fullRound <= io_input_payload_delay_66_fullRound;
    io_input_payload_delay_67_partialRound <= io_input_payload_delay_66_partialRound;
    io_input_payload_delay_67_stateIndex <= io_input_payload_delay_66_stateIndex;
    io_input_payload_delay_67_stateSize <= io_input_payload_delay_66_stateSize;
    io_input_payload_delay_67_stateID <= io_input_payload_delay_66_stateID;
    io_input_payload_delay_67_stateElements_0 <= io_input_payload_delay_66_stateElements_0;
    io_input_payload_delay_67_stateElements_1 <= io_input_payload_delay_66_stateElements_1;
    io_input_payload_delay_67_stateElements_2 <= io_input_payload_delay_66_stateElements_2;
    io_input_payload_delay_67_stateElements_3 <= io_input_payload_delay_66_stateElements_3;
    io_input_payload_delay_67_stateElements_4 <= io_input_payload_delay_66_stateElements_4;
    io_input_payload_delay_67_stateElements_5 <= io_input_payload_delay_66_stateElements_5;
    io_input_payload_delay_67_stateElements_6 <= io_input_payload_delay_66_stateElements_6;
    io_input_payload_delay_67_stateElements_7 <= io_input_payload_delay_66_stateElements_7;
    io_input_payload_delay_67_stateElements_8 <= io_input_payload_delay_66_stateElements_8;
    io_input_payload_delay_67_stateElements_9 <= io_input_payload_delay_66_stateElements_9;
    io_input_payload_delay_67_stateElements_10 <= io_input_payload_delay_66_stateElements_10;
    io_input_payload_delay_67_stateElement <= io_input_payload_delay_66_stateElement;
    io_input_payload_delay_68_isFull <= io_input_payload_delay_67_isFull;
    io_input_payload_delay_68_fullRound <= io_input_payload_delay_67_fullRound;
    io_input_payload_delay_68_partialRound <= io_input_payload_delay_67_partialRound;
    io_input_payload_delay_68_stateIndex <= io_input_payload_delay_67_stateIndex;
    io_input_payload_delay_68_stateSize <= io_input_payload_delay_67_stateSize;
    io_input_payload_delay_68_stateID <= io_input_payload_delay_67_stateID;
    io_input_payload_delay_68_stateElements_0 <= io_input_payload_delay_67_stateElements_0;
    io_input_payload_delay_68_stateElements_1 <= io_input_payload_delay_67_stateElements_1;
    io_input_payload_delay_68_stateElements_2 <= io_input_payload_delay_67_stateElements_2;
    io_input_payload_delay_68_stateElements_3 <= io_input_payload_delay_67_stateElements_3;
    io_input_payload_delay_68_stateElements_4 <= io_input_payload_delay_67_stateElements_4;
    io_input_payload_delay_68_stateElements_5 <= io_input_payload_delay_67_stateElements_5;
    io_input_payload_delay_68_stateElements_6 <= io_input_payload_delay_67_stateElements_6;
    io_input_payload_delay_68_stateElements_7 <= io_input_payload_delay_67_stateElements_7;
    io_input_payload_delay_68_stateElements_8 <= io_input_payload_delay_67_stateElements_8;
    io_input_payload_delay_68_stateElements_9 <= io_input_payload_delay_67_stateElements_9;
    io_input_payload_delay_68_stateElements_10 <= io_input_payload_delay_67_stateElements_10;
    io_input_payload_delay_68_stateElement <= io_input_payload_delay_67_stateElement;
    io_input_payload_delay_69_isFull <= io_input_payload_delay_68_isFull;
    io_input_payload_delay_69_fullRound <= io_input_payload_delay_68_fullRound;
    io_input_payload_delay_69_partialRound <= io_input_payload_delay_68_partialRound;
    io_input_payload_delay_69_stateIndex <= io_input_payload_delay_68_stateIndex;
    io_input_payload_delay_69_stateSize <= io_input_payload_delay_68_stateSize;
    io_input_payload_delay_69_stateID <= io_input_payload_delay_68_stateID;
    io_input_payload_delay_69_stateElements_0 <= io_input_payload_delay_68_stateElements_0;
    io_input_payload_delay_69_stateElements_1 <= io_input_payload_delay_68_stateElements_1;
    io_input_payload_delay_69_stateElements_2 <= io_input_payload_delay_68_stateElements_2;
    io_input_payload_delay_69_stateElements_3 <= io_input_payload_delay_68_stateElements_3;
    io_input_payload_delay_69_stateElements_4 <= io_input_payload_delay_68_stateElements_4;
    io_input_payload_delay_69_stateElements_5 <= io_input_payload_delay_68_stateElements_5;
    io_input_payload_delay_69_stateElements_6 <= io_input_payload_delay_68_stateElements_6;
    io_input_payload_delay_69_stateElements_7 <= io_input_payload_delay_68_stateElements_7;
    io_input_payload_delay_69_stateElements_8 <= io_input_payload_delay_68_stateElements_8;
    io_input_payload_delay_69_stateElements_9 <= io_input_payload_delay_68_stateElements_9;
    io_input_payload_delay_69_stateElements_10 <= io_input_payload_delay_68_stateElements_10;
    io_input_payload_delay_69_stateElement <= io_input_payload_delay_68_stateElement;
    io_input_payload_delay_70_isFull <= io_input_payload_delay_69_isFull;
    io_input_payload_delay_70_fullRound <= io_input_payload_delay_69_fullRound;
    io_input_payload_delay_70_partialRound <= io_input_payload_delay_69_partialRound;
    io_input_payload_delay_70_stateIndex <= io_input_payload_delay_69_stateIndex;
    io_input_payload_delay_70_stateSize <= io_input_payload_delay_69_stateSize;
    io_input_payload_delay_70_stateID <= io_input_payload_delay_69_stateID;
    io_input_payload_delay_70_stateElements_0 <= io_input_payload_delay_69_stateElements_0;
    io_input_payload_delay_70_stateElements_1 <= io_input_payload_delay_69_stateElements_1;
    io_input_payload_delay_70_stateElements_2 <= io_input_payload_delay_69_stateElements_2;
    io_input_payload_delay_70_stateElements_3 <= io_input_payload_delay_69_stateElements_3;
    io_input_payload_delay_70_stateElements_4 <= io_input_payload_delay_69_stateElements_4;
    io_input_payload_delay_70_stateElements_5 <= io_input_payload_delay_69_stateElements_5;
    io_input_payload_delay_70_stateElements_6 <= io_input_payload_delay_69_stateElements_6;
    io_input_payload_delay_70_stateElements_7 <= io_input_payload_delay_69_stateElements_7;
    io_input_payload_delay_70_stateElements_8 <= io_input_payload_delay_69_stateElements_8;
    io_input_payload_delay_70_stateElements_9 <= io_input_payload_delay_69_stateElements_9;
    io_input_payload_delay_70_stateElements_10 <= io_input_payload_delay_69_stateElements_10;
    io_input_payload_delay_70_stateElement <= io_input_payload_delay_69_stateElement;
    io_input_payload_delay_71_isFull <= io_input_payload_delay_70_isFull;
    io_input_payload_delay_71_fullRound <= io_input_payload_delay_70_fullRound;
    io_input_payload_delay_71_partialRound <= io_input_payload_delay_70_partialRound;
    io_input_payload_delay_71_stateIndex <= io_input_payload_delay_70_stateIndex;
    io_input_payload_delay_71_stateSize <= io_input_payload_delay_70_stateSize;
    io_input_payload_delay_71_stateID <= io_input_payload_delay_70_stateID;
    io_input_payload_delay_71_stateElements_0 <= io_input_payload_delay_70_stateElements_0;
    io_input_payload_delay_71_stateElements_1 <= io_input_payload_delay_70_stateElements_1;
    io_input_payload_delay_71_stateElements_2 <= io_input_payload_delay_70_stateElements_2;
    io_input_payload_delay_71_stateElements_3 <= io_input_payload_delay_70_stateElements_3;
    io_input_payload_delay_71_stateElements_4 <= io_input_payload_delay_70_stateElements_4;
    io_input_payload_delay_71_stateElements_5 <= io_input_payload_delay_70_stateElements_5;
    io_input_payload_delay_71_stateElements_6 <= io_input_payload_delay_70_stateElements_6;
    io_input_payload_delay_71_stateElements_7 <= io_input_payload_delay_70_stateElements_7;
    io_input_payload_delay_71_stateElements_8 <= io_input_payload_delay_70_stateElements_8;
    io_input_payload_delay_71_stateElements_9 <= io_input_payload_delay_70_stateElements_9;
    io_input_payload_delay_71_stateElements_10 <= io_input_payload_delay_70_stateElements_10;
    io_input_payload_delay_71_stateElement <= io_input_payload_delay_70_stateElement;
    io_input_payload_delay_72_isFull <= io_input_payload_delay_71_isFull;
    io_input_payload_delay_72_fullRound <= io_input_payload_delay_71_fullRound;
    io_input_payload_delay_72_partialRound <= io_input_payload_delay_71_partialRound;
    io_input_payload_delay_72_stateIndex <= io_input_payload_delay_71_stateIndex;
    io_input_payload_delay_72_stateSize <= io_input_payload_delay_71_stateSize;
    io_input_payload_delay_72_stateID <= io_input_payload_delay_71_stateID;
    io_input_payload_delay_72_stateElements_0 <= io_input_payload_delay_71_stateElements_0;
    io_input_payload_delay_72_stateElements_1 <= io_input_payload_delay_71_stateElements_1;
    io_input_payload_delay_72_stateElements_2 <= io_input_payload_delay_71_stateElements_2;
    io_input_payload_delay_72_stateElements_3 <= io_input_payload_delay_71_stateElements_3;
    io_input_payload_delay_72_stateElements_4 <= io_input_payload_delay_71_stateElements_4;
    io_input_payload_delay_72_stateElements_5 <= io_input_payload_delay_71_stateElements_5;
    io_input_payload_delay_72_stateElements_6 <= io_input_payload_delay_71_stateElements_6;
    io_input_payload_delay_72_stateElements_7 <= io_input_payload_delay_71_stateElements_7;
    io_input_payload_delay_72_stateElements_8 <= io_input_payload_delay_71_stateElements_8;
    io_input_payload_delay_72_stateElements_9 <= io_input_payload_delay_71_stateElements_9;
    io_input_payload_delay_72_stateElements_10 <= io_input_payload_delay_71_stateElements_10;
    io_input_payload_delay_72_stateElement <= io_input_payload_delay_71_stateElement;
    io_input_payload_delay_73_isFull <= io_input_payload_delay_72_isFull;
    io_input_payload_delay_73_fullRound <= io_input_payload_delay_72_fullRound;
    io_input_payload_delay_73_partialRound <= io_input_payload_delay_72_partialRound;
    io_input_payload_delay_73_stateIndex <= io_input_payload_delay_72_stateIndex;
    io_input_payload_delay_73_stateSize <= io_input_payload_delay_72_stateSize;
    io_input_payload_delay_73_stateID <= io_input_payload_delay_72_stateID;
    io_input_payload_delay_73_stateElements_0 <= io_input_payload_delay_72_stateElements_0;
    io_input_payload_delay_73_stateElements_1 <= io_input_payload_delay_72_stateElements_1;
    io_input_payload_delay_73_stateElements_2 <= io_input_payload_delay_72_stateElements_2;
    io_input_payload_delay_73_stateElements_3 <= io_input_payload_delay_72_stateElements_3;
    io_input_payload_delay_73_stateElements_4 <= io_input_payload_delay_72_stateElements_4;
    io_input_payload_delay_73_stateElements_5 <= io_input_payload_delay_72_stateElements_5;
    io_input_payload_delay_73_stateElements_6 <= io_input_payload_delay_72_stateElements_6;
    io_input_payload_delay_73_stateElements_7 <= io_input_payload_delay_72_stateElements_7;
    io_input_payload_delay_73_stateElements_8 <= io_input_payload_delay_72_stateElements_8;
    io_input_payload_delay_73_stateElements_9 <= io_input_payload_delay_72_stateElements_9;
    io_input_payload_delay_73_stateElements_10 <= io_input_payload_delay_72_stateElements_10;
    io_input_payload_delay_73_stateElement <= io_input_payload_delay_72_stateElement;
    io_input_payload_delay_74_isFull <= io_input_payload_delay_73_isFull;
    io_input_payload_delay_74_fullRound <= io_input_payload_delay_73_fullRound;
    io_input_payload_delay_74_partialRound <= io_input_payload_delay_73_partialRound;
    io_input_payload_delay_74_stateIndex <= io_input_payload_delay_73_stateIndex;
    io_input_payload_delay_74_stateSize <= io_input_payload_delay_73_stateSize;
    io_input_payload_delay_74_stateID <= io_input_payload_delay_73_stateID;
    io_input_payload_delay_74_stateElements_0 <= io_input_payload_delay_73_stateElements_0;
    io_input_payload_delay_74_stateElements_1 <= io_input_payload_delay_73_stateElements_1;
    io_input_payload_delay_74_stateElements_2 <= io_input_payload_delay_73_stateElements_2;
    io_input_payload_delay_74_stateElements_3 <= io_input_payload_delay_73_stateElements_3;
    io_input_payload_delay_74_stateElements_4 <= io_input_payload_delay_73_stateElements_4;
    io_input_payload_delay_74_stateElements_5 <= io_input_payload_delay_73_stateElements_5;
    io_input_payload_delay_74_stateElements_6 <= io_input_payload_delay_73_stateElements_6;
    io_input_payload_delay_74_stateElements_7 <= io_input_payload_delay_73_stateElements_7;
    io_input_payload_delay_74_stateElements_8 <= io_input_payload_delay_73_stateElements_8;
    io_input_payload_delay_74_stateElements_9 <= io_input_payload_delay_73_stateElements_9;
    io_input_payload_delay_74_stateElements_10 <= io_input_payload_delay_73_stateElements_10;
    io_input_payload_delay_74_stateElement <= io_input_payload_delay_73_stateElement;
    io_input_payload_delay_75_isFull <= io_input_payload_delay_74_isFull;
    io_input_payload_delay_75_fullRound <= io_input_payload_delay_74_fullRound;
    io_input_payload_delay_75_partialRound <= io_input_payload_delay_74_partialRound;
    io_input_payload_delay_75_stateIndex <= io_input_payload_delay_74_stateIndex;
    io_input_payload_delay_75_stateSize <= io_input_payload_delay_74_stateSize;
    io_input_payload_delay_75_stateID <= io_input_payload_delay_74_stateID;
    io_input_payload_delay_75_stateElements_0 <= io_input_payload_delay_74_stateElements_0;
    io_input_payload_delay_75_stateElements_1 <= io_input_payload_delay_74_stateElements_1;
    io_input_payload_delay_75_stateElements_2 <= io_input_payload_delay_74_stateElements_2;
    io_input_payload_delay_75_stateElements_3 <= io_input_payload_delay_74_stateElements_3;
    io_input_payload_delay_75_stateElements_4 <= io_input_payload_delay_74_stateElements_4;
    io_input_payload_delay_75_stateElements_5 <= io_input_payload_delay_74_stateElements_5;
    io_input_payload_delay_75_stateElements_6 <= io_input_payload_delay_74_stateElements_6;
    io_input_payload_delay_75_stateElements_7 <= io_input_payload_delay_74_stateElements_7;
    io_input_payload_delay_75_stateElements_8 <= io_input_payload_delay_74_stateElements_8;
    io_input_payload_delay_75_stateElements_9 <= io_input_payload_delay_74_stateElements_9;
    io_input_payload_delay_75_stateElements_10 <= io_input_payload_delay_74_stateElements_10;
    io_input_payload_delay_75_stateElement <= io_input_payload_delay_74_stateElement;
    io_input_payload_delay_76_isFull <= io_input_payload_delay_75_isFull;
    io_input_payload_delay_76_fullRound <= io_input_payload_delay_75_fullRound;
    io_input_payload_delay_76_partialRound <= io_input_payload_delay_75_partialRound;
    io_input_payload_delay_76_stateIndex <= io_input_payload_delay_75_stateIndex;
    io_input_payload_delay_76_stateSize <= io_input_payload_delay_75_stateSize;
    io_input_payload_delay_76_stateID <= io_input_payload_delay_75_stateID;
    io_input_payload_delay_76_stateElements_0 <= io_input_payload_delay_75_stateElements_0;
    io_input_payload_delay_76_stateElements_1 <= io_input_payload_delay_75_stateElements_1;
    io_input_payload_delay_76_stateElements_2 <= io_input_payload_delay_75_stateElements_2;
    io_input_payload_delay_76_stateElements_3 <= io_input_payload_delay_75_stateElements_3;
    io_input_payload_delay_76_stateElements_4 <= io_input_payload_delay_75_stateElements_4;
    io_input_payload_delay_76_stateElements_5 <= io_input_payload_delay_75_stateElements_5;
    io_input_payload_delay_76_stateElements_6 <= io_input_payload_delay_75_stateElements_6;
    io_input_payload_delay_76_stateElements_7 <= io_input_payload_delay_75_stateElements_7;
    io_input_payload_delay_76_stateElements_8 <= io_input_payload_delay_75_stateElements_8;
    io_input_payload_delay_76_stateElements_9 <= io_input_payload_delay_75_stateElements_9;
    io_input_payload_delay_76_stateElements_10 <= io_input_payload_delay_75_stateElements_10;
    io_input_payload_delay_76_stateElement <= io_input_payload_delay_75_stateElement;
    io_input_payload_delay_77_isFull <= io_input_payload_delay_76_isFull;
    io_input_payload_delay_77_fullRound <= io_input_payload_delay_76_fullRound;
    io_input_payload_delay_77_partialRound <= io_input_payload_delay_76_partialRound;
    io_input_payload_delay_77_stateIndex <= io_input_payload_delay_76_stateIndex;
    io_input_payload_delay_77_stateSize <= io_input_payload_delay_76_stateSize;
    io_input_payload_delay_77_stateID <= io_input_payload_delay_76_stateID;
    io_input_payload_delay_77_stateElements_0 <= io_input_payload_delay_76_stateElements_0;
    io_input_payload_delay_77_stateElements_1 <= io_input_payload_delay_76_stateElements_1;
    io_input_payload_delay_77_stateElements_2 <= io_input_payload_delay_76_stateElements_2;
    io_input_payload_delay_77_stateElements_3 <= io_input_payload_delay_76_stateElements_3;
    io_input_payload_delay_77_stateElements_4 <= io_input_payload_delay_76_stateElements_4;
    io_input_payload_delay_77_stateElements_5 <= io_input_payload_delay_76_stateElements_5;
    io_input_payload_delay_77_stateElements_6 <= io_input_payload_delay_76_stateElements_6;
    io_input_payload_delay_77_stateElements_7 <= io_input_payload_delay_76_stateElements_7;
    io_input_payload_delay_77_stateElements_8 <= io_input_payload_delay_76_stateElements_8;
    io_input_payload_delay_77_stateElements_9 <= io_input_payload_delay_76_stateElements_9;
    io_input_payload_delay_77_stateElements_10 <= io_input_payload_delay_76_stateElements_10;
    io_input_payload_delay_77_stateElement <= io_input_payload_delay_76_stateElement;
    io_input_payload_delay_78_isFull <= io_input_payload_delay_77_isFull;
    io_input_payload_delay_78_fullRound <= io_input_payload_delay_77_fullRound;
    io_input_payload_delay_78_partialRound <= io_input_payload_delay_77_partialRound;
    io_input_payload_delay_78_stateIndex <= io_input_payload_delay_77_stateIndex;
    io_input_payload_delay_78_stateSize <= io_input_payload_delay_77_stateSize;
    io_input_payload_delay_78_stateID <= io_input_payload_delay_77_stateID;
    io_input_payload_delay_78_stateElements_0 <= io_input_payload_delay_77_stateElements_0;
    io_input_payload_delay_78_stateElements_1 <= io_input_payload_delay_77_stateElements_1;
    io_input_payload_delay_78_stateElements_2 <= io_input_payload_delay_77_stateElements_2;
    io_input_payload_delay_78_stateElements_3 <= io_input_payload_delay_77_stateElements_3;
    io_input_payload_delay_78_stateElements_4 <= io_input_payload_delay_77_stateElements_4;
    io_input_payload_delay_78_stateElements_5 <= io_input_payload_delay_77_stateElements_5;
    io_input_payload_delay_78_stateElements_6 <= io_input_payload_delay_77_stateElements_6;
    io_input_payload_delay_78_stateElements_7 <= io_input_payload_delay_77_stateElements_7;
    io_input_payload_delay_78_stateElements_8 <= io_input_payload_delay_77_stateElements_8;
    io_input_payload_delay_78_stateElements_9 <= io_input_payload_delay_77_stateElements_9;
    io_input_payload_delay_78_stateElements_10 <= io_input_payload_delay_77_stateElements_10;
    io_input_payload_delay_78_stateElement <= io_input_payload_delay_77_stateElement;
    io_input_payload_delay_79_isFull <= io_input_payload_delay_78_isFull;
    io_input_payload_delay_79_fullRound <= io_input_payload_delay_78_fullRound;
    io_input_payload_delay_79_partialRound <= io_input_payload_delay_78_partialRound;
    io_input_payload_delay_79_stateIndex <= io_input_payload_delay_78_stateIndex;
    io_input_payload_delay_79_stateSize <= io_input_payload_delay_78_stateSize;
    io_input_payload_delay_79_stateID <= io_input_payload_delay_78_stateID;
    io_input_payload_delay_79_stateElements_0 <= io_input_payload_delay_78_stateElements_0;
    io_input_payload_delay_79_stateElements_1 <= io_input_payload_delay_78_stateElements_1;
    io_input_payload_delay_79_stateElements_2 <= io_input_payload_delay_78_stateElements_2;
    io_input_payload_delay_79_stateElements_3 <= io_input_payload_delay_78_stateElements_3;
    io_input_payload_delay_79_stateElements_4 <= io_input_payload_delay_78_stateElements_4;
    io_input_payload_delay_79_stateElements_5 <= io_input_payload_delay_78_stateElements_5;
    io_input_payload_delay_79_stateElements_6 <= io_input_payload_delay_78_stateElements_6;
    io_input_payload_delay_79_stateElements_7 <= io_input_payload_delay_78_stateElements_7;
    io_input_payload_delay_79_stateElements_8 <= io_input_payload_delay_78_stateElements_8;
    io_input_payload_delay_79_stateElements_9 <= io_input_payload_delay_78_stateElements_9;
    io_input_payload_delay_79_stateElements_10 <= io_input_payload_delay_78_stateElements_10;
    io_input_payload_delay_79_stateElement <= io_input_payload_delay_78_stateElement;
    io_input_payload_delay_80_isFull <= io_input_payload_delay_79_isFull;
    io_input_payload_delay_80_fullRound <= io_input_payload_delay_79_fullRound;
    io_input_payload_delay_80_partialRound <= io_input_payload_delay_79_partialRound;
    io_input_payload_delay_80_stateIndex <= io_input_payload_delay_79_stateIndex;
    io_input_payload_delay_80_stateSize <= io_input_payload_delay_79_stateSize;
    io_input_payload_delay_80_stateID <= io_input_payload_delay_79_stateID;
    io_input_payload_delay_80_stateElements_0 <= io_input_payload_delay_79_stateElements_0;
    io_input_payload_delay_80_stateElements_1 <= io_input_payload_delay_79_stateElements_1;
    io_input_payload_delay_80_stateElements_2 <= io_input_payload_delay_79_stateElements_2;
    io_input_payload_delay_80_stateElements_3 <= io_input_payload_delay_79_stateElements_3;
    io_input_payload_delay_80_stateElements_4 <= io_input_payload_delay_79_stateElements_4;
    io_input_payload_delay_80_stateElements_5 <= io_input_payload_delay_79_stateElements_5;
    io_input_payload_delay_80_stateElements_6 <= io_input_payload_delay_79_stateElements_6;
    io_input_payload_delay_80_stateElements_7 <= io_input_payload_delay_79_stateElements_7;
    io_input_payload_delay_80_stateElements_8 <= io_input_payload_delay_79_stateElements_8;
    io_input_payload_delay_80_stateElements_9 <= io_input_payload_delay_79_stateElements_9;
    io_input_payload_delay_80_stateElements_10 <= io_input_payload_delay_79_stateElements_10;
    io_input_payload_delay_80_stateElement <= io_input_payload_delay_79_stateElement;
    io_input_payload_delay_81_isFull <= io_input_payload_delay_80_isFull;
    io_input_payload_delay_81_fullRound <= io_input_payload_delay_80_fullRound;
    io_input_payload_delay_81_partialRound <= io_input_payload_delay_80_partialRound;
    io_input_payload_delay_81_stateIndex <= io_input_payload_delay_80_stateIndex;
    io_input_payload_delay_81_stateSize <= io_input_payload_delay_80_stateSize;
    io_input_payload_delay_81_stateID <= io_input_payload_delay_80_stateID;
    io_input_payload_delay_81_stateElements_0 <= io_input_payload_delay_80_stateElements_0;
    io_input_payload_delay_81_stateElements_1 <= io_input_payload_delay_80_stateElements_1;
    io_input_payload_delay_81_stateElements_2 <= io_input_payload_delay_80_stateElements_2;
    io_input_payload_delay_81_stateElements_3 <= io_input_payload_delay_80_stateElements_3;
    io_input_payload_delay_81_stateElements_4 <= io_input_payload_delay_80_stateElements_4;
    io_input_payload_delay_81_stateElements_5 <= io_input_payload_delay_80_stateElements_5;
    io_input_payload_delay_81_stateElements_6 <= io_input_payload_delay_80_stateElements_6;
    io_input_payload_delay_81_stateElements_7 <= io_input_payload_delay_80_stateElements_7;
    io_input_payload_delay_81_stateElements_8 <= io_input_payload_delay_80_stateElements_8;
    io_input_payload_delay_81_stateElements_9 <= io_input_payload_delay_80_stateElements_9;
    io_input_payload_delay_81_stateElements_10 <= io_input_payload_delay_80_stateElements_10;
    io_input_payload_delay_81_stateElement <= io_input_payload_delay_80_stateElement;
    io_input_payload_delay_82_isFull <= io_input_payload_delay_81_isFull;
    io_input_payload_delay_82_fullRound <= io_input_payload_delay_81_fullRound;
    io_input_payload_delay_82_partialRound <= io_input_payload_delay_81_partialRound;
    io_input_payload_delay_82_stateIndex <= io_input_payload_delay_81_stateIndex;
    io_input_payload_delay_82_stateSize <= io_input_payload_delay_81_stateSize;
    io_input_payload_delay_82_stateID <= io_input_payload_delay_81_stateID;
    io_input_payload_delay_82_stateElements_0 <= io_input_payload_delay_81_stateElements_0;
    io_input_payload_delay_82_stateElements_1 <= io_input_payload_delay_81_stateElements_1;
    io_input_payload_delay_82_stateElements_2 <= io_input_payload_delay_81_stateElements_2;
    io_input_payload_delay_82_stateElements_3 <= io_input_payload_delay_81_stateElements_3;
    io_input_payload_delay_82_stateElements_4 <= io_input_payload_delay_81_stateElements_4;
    io_input_payload_delay_82_stateElements_5 <= io_input_payload_delay_81_stateElements_5;
    io_input_payload_delay_82_stateElements_6 <= io_input_payload_delay_81_stateElements_6;
    io_input_payload_delay_82_stateElements_7 <= io_input_payload_delay_81_stateElements_7;
    io_input_payload_delay_82_stateElements_8 <= io_input_payload_delay_81_stateElements_8;
    io_input_payload_delay_82_stateElements_9 <= io_input_payload_delay_81_stateElements_9;
    io_input_payload_delay_82_stateElements_10 <= io_input_payload_delay_81_stateElements_10;
    io_input_payload_delay_82_stateElement <= io_input_payload_delay_81_stateElement;
    io_input_payload_delay_83_isFull <= io_input_payload_delay_82_isFull;
    io_input_payload_delay_83_fullRound <= io_input_payload_delay_82_fullRound;
    io_input_payload_delay_83_partialRound <= io_input_payload_delay_82_partialRound;
    io_input_payload_delay_83_stateIndex <= io_input_payload_delay_82_stateIndex;
    io_input_payload_delay_83_stateSize <= io_input_payload_delay_82_stateSize;
    io_input_payload_delay_83_stateID <= io_input_payload_delay_82_stateID;
    io_input_payload_delay_83_stateElements_0 <= io_input_payload_delay_82_stateElements_0;
    io_input_payload_delay_83_stateElements_1 <= io_input_payload_delay_82_stateElements_1;
    io_input_payload_delay_83_stateElements_2 <= io_input_payload_delay_82_stateElements_2;
    io_input_payload_delay_83_stateElements_3 <= io_input_payload_delay_82_stateElements_3;
    io_input_payload_delay_83_stateElements_4 <= io_input_payload_delay_82_stateElements_4;
    io_input_payload_delay_83_stateElements_5 <= io_input_payload_delay_82_stateElements_5;
    io_input_payload_delay_83_stateElements_6 <= io_input_payload_delay_82_stateElements_6;
    io_input_payload_delay_83_stateElements_7 <= io_input_payload_delay_82_stateElements_7;
    io_input_payload_delay_83_stateElements_8 <= io_input_payload_delay_82_stateElements_8;
    io_input_payload_delay_83_stateElements_9 <= io_input_payload_delay_82_stateElements_9;
    io_input_payload_delay_83_stateElements_10 <= io_input_payload_delay_82_stateElements_10;
    io_input_payload_delay_83_stateElement <= io_input_payload_delay_82_stateElement;
    io_input_payload_delay_84_isFull <= io_input_payload_delay_83_isFull;
    io_input_payload_delay_84_fullRound <= io_input_payload_delay_83_fullRound;
    io_input_payload_delay_84_partialRound <= io_input_payload_delay_83_partialRound;
    io_input_payload_delay_84_stateIndex <= io_input_payload_delay_83_stateIndex;
    io_input_payload_delay_84_stateSize <= io_input_payload_delay_83_stateSize;
    io_input_payload_delay_84_stateID <= io_input_payload_delay_83_stateID;
    io_input_payload_delay_84_stateElements_0 <= io_input_payload_delay_83_stateElements_0;
    io_input_payload_delay_84_stateElements_1 <= io_input_payload_delay_83_stateElements_1;
    io_input_payload_delay_84_stateElements_2 <= io_input_payload_delay_83_stateElements_2;
    io_input_payload_delay_84_stateElements_3 <= io_input_payload_delay_83_stateElements_3;
    io_input_payload_delay_84_stateElements_4 <= io_input_payload_delay_83_stateElements_4;
    io_input_payload_delay_84_stateElements_5 <= io_input_payload_delay_83_stateElements_5;
    io_input_payload_delay_84_stateElements_6 <= io_input_payload_delay_83_stateElements_6;
    io_input_payload_delay_84_stateElements_7 <= io_input_payload_delay_83_stateElements_7;
    io_input_payload_delay_84_stateElements_8 <= io_input_payload_delay_83_stateElements_8;
    io_input_payload_delay_84_stateElements_9 <= io_input_payload_delay_83_stateElements_9;
    io_input_payload_delay_84_stateElements_10 <= io_input_payload_delay_83_stateElements_10;
    io_input_payload_delay_84_stateElement <= io_input_payload_delay_83_stateElement;
    io_input_payload_delay_85_isFull <= io_input_payload_delay_84_isFull;
    io_input_payload_delay_85_fullRound <= io_input_payload_delay_84_fullRound;
    io_input_payload_delay_85_partialRound <= io_input_payload_delay_84_partialRound;
    io_input_payload_delay_85_stateIndex <= io_input_payload_delay_84_stateIndex;
    io_input_payload_delay_85_stateSize <= io_input_payload_delay_84_stateSize;
    io_input_payload_delay_85_stateID <= io_input_payload_delay_84_stateID;
    io_input_payload_delay_85_stateElements_0 <= io_input_payload_delay_84_stateElements_0;
    io_input_payload_delay_85_stateElements_1 <= io_input_payload_delay_84_stateElements_1;
    io_input_payload_delay_85_stateElements_2 <= io_input_payload_delay_84_stateElements_2;
    io_input_payload_delay_85_stateElements_3 <= io_input_payload_delay_84_stateElements_3;
    io_input_payload_delay_85_stateElements_4 <= io_input_payload_delay_84_stateElements_4;
    io_input_payload_delay_85_stateElements_5 <= io_input_payload_delay_84_stateElements_5;
    io_input_payload_delay_85_stateElements_6 <= io_input_payload_delay_84_stateElements_6;
    io_input_payload_delay_85_stateElements_7 <= io_input_payload_delay_84_stateElements_7;
    io_input_payload_delay_85_stateElements_8 <= io_input_payload_delay_84_stateElements_8;
    io_input_payload_delay_85_stateElements_9 <= io_input_payload_delay_84_stateElements_9;
    io_input_payload_delay_85_stateElements_10 <= io_input_payload_delay_84_stateElements_10;
    io_input_payload_delay_85_stateElement <= io_input_payload_delay_84_stateElement;
    io_input_payload_delay_86_isFull <= io_input_payload_delay_85_isFull;
    io_input_payload_delay_86_fullRound <= io_input_payload_delay_85_fullRound;
    io_input_payload_delay_86_partialRound <= io_input_payload_delay_85_partialRound;
    io_input_payload_delay_86_stateIndex <= io_input_payload_delay_85_stateIndex;
    io_input_payload_delay_86_stateSize <= io_input_payload_delay_85_stateSize;
    io_input_payload_delay_86_stateID <= io_input_payload_delay_85_stateID;
    io_input_payload_delay_86_stateElements_0 <= io_input_payload_delay_85_stateElements_0;
    io_input_payload_delay_86_stateElements_1 <= io_input_payload_delay_85_stateElements_1;
    io_input_payload_delay_86_stateElements_2 <= io_input_payload_delay_85_stateElements_2;
    io_input_payload_delay_86_stateElements_3 <= io_input_payload_delay_85_stateElements_3;
    io_input_payload_delay_86_stateElements_4 <= io_input_payload_delay_85_stateElements_4;
    io_input_payload_delay_86_stateElements_5 <= io_input_payload_delay_85_stateElements_5;
    io_input_payload_delay_86_stateElements_6 <= io_input_payload_delay_85_stateElements_6;
    io_input_payload_delay_86_stateElements_7 <= io_input_payload_delay_85_stateElements_7;
    io_input_payload_delay_86_stateElements_8 <= io_input_payload_delay_85_stateElements_8;
    io_input_payload_delay_86_stateElements_9 <= io_input_payload_delay_85_stateElements_9;
    io_input_payload_delay_86_stateElements_10 <= io_input_payload_delay_85_stateElements_10;
    io_input_payload_delay_86_stateElement <= io_input_payload_delay_85_stateElement;
    io_input_payload_delay_87_isFull <= io_input_payload_delay_86_isFull;
    io_input_payload_delay_87_fullRound <= io_input_payload_delay_86_fullRound;
    io_input_payload_delay_87_partialRound <= io_input_payload_delay_86_partialRound;
    io_input_payload_delay_87_stateIndex <= io_input_payload_delay_86_stateIndex;
    io_input_payload_delay_87_stateSize <= io_input_payload_delay_86_stateSize;
    io_input_payload_delay_87_stateID <= io_input_payload_delay_86_stateID;
    io_input_payload_delay_87_stateElements_0 <= io_input_payload_delay_86_stateElements_0;
    io_input_payload_delay_87_stateElements_1 <= io_input_payload_delay_86_stateElements_1;
    io_input_payload_delay_87_stateElements_2 <= io_input_payload_delay_86_stateElements_2;
    io_input_payload_delay_87_stateElements_3 <= io_input_payload_delay_86_stateElements_3;
    io_input_payload_delay_87_stateElements_4 <= io_input_payload_delay_86_stateElements_4;
    io_input_payload_delay_87_stateElements_5 <= io_input_payload_delay_86_stateElements_5;
    io_input_payload_delay_87_stateElements_6 <= io_input_payload_delay_86_stateElements_6;
    io_input_payload_delay_87_stateElements_7 <= io_input_payload_delay_86_stateElements_7;
    io_input_payload_delay_87_stateElements_8 <= io_input_payload_delay_86_stateElements_8;
    io_input_payload_delay_87_stateElements_9 <= io_input_payload_delay_86_stateElements_9;
    io_input_payload_delay_87_stateElements_10 <= io_input_payload_delay_86_stateElements_10;
    io_input_payload_delay_87_stateElement <= io_input_payload_delay_86_stateElement;
    io_input_payload_delay_88_isFull <= io_input_payload_delay_87_isFull;
    io_input_payload_delay_88_fullRound <= io_input_payload_delay_87_fullRound;
    io_input_payload_delay_88_partialRound <= io_input_payload_delay_87_partialRound;
    io_input_payload_delay_88_stateIndex <= io_input_payload_delay_87_stateIndex;
    io_input_payload_delay_88_stateSize <= io_input_payload_delay_87_stateSize;
    io_input_payload_delay_88_stateID <= io_input_payload_delay_87_stateID;
    io_input_payload_delay_88_stateElements_0 <= io_input_payload_delay_87_stateElements_0;
    io_input_payload_delay_88_stateElements_1 <= io_input_payload_delay_87_stateElements_1;
    io_input_payload_delay_88_stateElements_2 <= io_input_payload_delay_87_stateElements_2;
    io_input_payload_delay_88_stateElements_3 <= io_input_payload_delay_87_stateElements_3;
    io_input_payload_delay_88_stateElements_4 <= io_input_payload_delay_87_stateElements_4;
    io_input_payload_delay_88_stateElements_5 <= io_input_payload_delay_87_stateElements_5;
    io_input_payload_delay_88_stateElements_6 <= io_input_payload_delay_87_stateElements_6;
    io_input_payload_delay_88_stateElements_7 <= io_input_payload_delay_87_stateElements_7;
    io_input_payload_delay_88_stateElements_8 <= io_input_payload_delay_87_stateElements_8;
    io_input_payload_delay_88_stateElements_9 <= io_input_payload_delay_87_stateElements_9;
    io_input_payload_delay_88_stateElements_10 <= io_input_payload_delay_87_stateElements_10;
    io_input_payload_delay_88_stateElement <= io_input_payload_delay_87_stateElement;
    io_input_payload_delay_89_isFull <= io_input_payload_delay_88_isFull;
    io_input_payload_delay_89_fullRound <= io_input_payload_delay_88_fullRound;
    io_input_payload_delay_89_partialRound <= io_input_payload_delay_88_partialRound;
    io_input_payload_delay_89_stateIndex <= io_input_payload_delay_88_stateIndex;
    io_input_payload_delay_89_stateSize <= io_input_payload_delay_88_stateSize;
    io_input_payload_delay_89_stateID <= io_input_payload_delay_88_stateID;
    io_input_payload_delay_89_stateElements_0 <= io_input_payload_delay_88_stateElements_0;
    io_input_payload_delay_89_stateElements_1 <= io_input_payload_delay_88_stateElements_1;
    io_input_payload_delay_89_stateElements_2 <= io_input_payload_delay_88_stateElements_2;
    io_input_payload_delay_89_stateElements_3 <= io_input_payload_delay_88_stateElements_3;
    io_input_payload_delay_89_stateElements_4 <= io_input_payload_delay_88_stateElements_4;
    io_input_payload_delay_89_stateElements_5 <= io_input_payload_delay_88_stateElements_5;
    io_input_payload_delay_89_stateElements_6 <= io_input_payload_delay_88_stateElements_6;
    io_input_payload_delay_89_stateElements_7 <= io_input_payload_delay_88_stateElements_7;
    io_input_payload_delay_89_stateElements_8 <= io_input_payload_delay_88_stateElements_8;
    io_input_payload_delay_89_stateElements_9 <= io_input_payload_delay_88_stateElements_9;
    io_input_payload_delay_89_stateElements_10 <= io_input_payload_delay_88_stateElements_10;
    io_input_payload_delay_89_stateElement <= io_input_payload_delay_88_stateElement;
    io_input_payload_delay_90_isFull <= io_input_payload_delay_89_isFull;
    io_input_payload_delay_90_fullRound <= io_input_payload_delay_89_fullRound;
    io_input_payload_delay_90_partialRound <= io_input_payload_delay_89_partialRound;
    io_input_payload_delay_90_stateIndex <= io_input_payload_delay_89_stateIndex;
    io_input_payload_delay_90_stateSize <= io_input_payload_delay_89_stateSize;
    io_input_payload_delay_90_stateID <= io_input_payload_delay_89_stateID;
    io_input_payload_delay_90_stateElements_0 <= io_input_payload_delay_89_stateElements_0;
    io_input_payload_delay_90_stateElements_1 <= io_input_payload_delay_89_stateElements_1;
    io_input_payload_delay_90_stateElements_2 <= io_input_payload_delay_89_stateElements_2;
    io_input_payload_delay_90_stateElements_3 <= io_input_payload_delay_89_stateElements_3;
    io_input_payload_delay_90_stateElements_4 <= io_input_payload_delay_89_stateElements_4;
    io_input_payload_delay_90_stateElements_5 <= io_input_payload_delay_89_stateElements_5;
    io_input_payload_delay_90_stateElements_6 <= io_input_payload_delay_89_stateElements_6;
    io_input_payload_delay_90_stateElements_7 <= io_input_payload_delay_89_stateElements_7;
    io_input_payload_delay_90_stateElements_8 <= io_input_payload_delay_89_stateElements_8;
    io_input_payload_delay_90_stateElements_9 <= io_input_payload_delay_89_stateElements_9;
    io_input_payload_delay_90_stateElements_10 <= io_input_payload_delay_89_stateElements_10;
    io_input_payload_delay_90_stateElement <= io_input_payload_delay_89_stateElement;
    io_input_payload_delay_91_isFull <= io_input_payload_delay_90_isFull;
    io_input_payload_delay_91_fullRound <= io_input_payload_delay_90_fullRound;
    io_input_payload_delay_91_partialRound <= io_input_payload_delay_90_partialRound;
    io_input_payload_delay_91_stateIndex <= io_input_payload_delay_90_stateIndex;
    io_input_payload_delay_91_stateSize <= io_input_payload_delay_90_stateSize;
    io_input_payload_delay_91_stateID <= io_input_payload_delay_90_stateID;
    io_input_payload_delay_91_stateElements_0 <= io_input_payload_delay_90_stateElements_0;
    io_input_payload_delay_91_stateElements_1 <= io_input_payload_delay_90_stateElements_1;
    io_input_payload_delay_91_stateElements_2 <= io_input_payload_delay_90_stateElements_2;
    io_input_payload_delay_91_stateElements_3 <= io_input_payload_delay_90_stateElements_3;
    io_input_payload_delay_91_stateElements_4 <= io_input_payload_delay_90_stateElements_4;
    io_input_payload_delay_91_stateElements_5 <= io_input_payload_delay_90_stateElements_5;
    io_input_payload_delay_91_stateElements_6 <= io_input_payload_delay_90_stateElements_6;
    io_input_payload_delay_91_stateElements_7 <= io_input_payload_delay_90_stateElements_7;
    io_input_payload_delay_91_stateElements_8 <= io_input_payload_delay_90_stateElements_8;
    io_input_payload_delay_91_stateElements_9 <= io_input_payload_delay_90_stateElements_9;
    io_input_payload_delay_91_stateElements_10 <= io_input_payload_delay_90_stateElements_10;
    io_input_payload_delay_91_stateElement <= io_input_payload_delay_90_stateElement;
    io_input_payload_delay_92_isFull <= io_input_payload_delay_91_isFull;
    io_input_payload_delay_92_fullRound <= io_input_payload_delay_91_fullRound;
    io_input_payload_delay_92_partialRound <= io_input_payload_delay_91_partialRound;
    io_input_payload_delay_92_stateIndex <= io_input_payload_delay_91_stateIndex;
    io_input_payload_delay_92_stateSize <= io_input_payload_delay_91_stateSize;
    io_input_payload_delay_92_stateID <= io_input_payload_delay_91_stateID;
    io_input_payload_delay_92_stateElements_0 <= io_input_payload_delay_91_stateElements_0;
    io_input_payload_delay_92_stateElements_1 <= io_input_payload_delay_91_stateElements_1;
    io_input_payload_delay_92_stateElements_2 <= io_input_payload_delay_91_stateElements_2;
    io_input_payload_delay_92_stateElements_3 <= io_input_payload_delay_91_stateElements_3;
    io_input_payload_delay_92_stateElements_4 <= io_input_payload_delay_91_stateElements_4;
    io_input_payload_delay_92_stateElements_5 <= io_input_payload_delay_91_stateElements_5;
    io_input_payload_delay_92_stateElements_6 <= io_input_payload_delay_91_stateElements_6;
    io_input_payload_delay_92_stateElements_7 <= io_input_payload_delay_91_stateElements_7;
    io_input_payload_delay_92_stateElements_8 <= io_input_payload_delay_91_stateElements_8;
    io_input_payload_delay_92_stateElements_9 <= io_input_payload_delay_91_stateElements_9;
    io_input_payload_delay_92_stateElements_10 <= io_input_payload_delay_91_stateElements_10;
    io_input_payload_delay_92_stateElement <= io_input_payload_delay_91_stateElement;
    io_input_payload_delay_93_isFull <= io_input_payload_delay_92_isFull;
    io_input_payload_delay_93_fullRound <= io_input_payload_delay_92_fullRound;
    io_input_payload_delay_93_partialRound <= io_input_payload_delay_92_partialRound;
    io_input_payload_delay_93_stateIndex <= io_input_payload_delay_92_stateIndex;
    io_input_payload_delay_93_stateSize <= io_input_payload_delay_92_stateSize;
    io_input_payload_delay_93_stateID <= io_input_payload_delay_92_stateID;
    io_input_payload_delay_93_stateElements_0 <= io_input_payload_delay_92_stateElements_0;
    io_input_payload_delay_93_stateElements_1 <= io_input_payload_delay_92_stateElements_1;
    io_input_payload_delay_93_stateElements_2 <= io_input_payload_delay_92_stateElements_2;
    io_input_payload_delay_93_stateElements_3 <= io_input_payload_delay_92_stateElements_3;
    io_input_payload_delay_93_stateElements_4 <= io_input_payload_delay_92_stateElements_4;
    io_input_payload_delay_93_stateElements_5 <= io_input_payload_delay_92_stateElements_5;
    io_input_payload_delay_93_stateElements_6 <= io_input_payload_delay_92_stateElements_6;
    io_input_payload_delay_93_stateElements_7 <= io_input_payload_delay_92_stateElements_7;
    io_input_payload_delay_93_stateElements_8 <= io_input_payload_delay_92_stateElements_8;
    io_input_payload_delay_93_stateElements_9 <= io_input_payload_delay_92_stateElements_9;
    io_input_payload_delay_93_stateElements_10 <= io_input_payload_delay_92_stateElements_10;
    io_input_payload_delay_93_stateElement <= io_input_payload_delay_92_stateElement;
    io_input_payload_delay_94_isFull <= io_input_payload_delay_93_isFull;
    io_input_payload_delay_94_fullRound <= io_input_payload_delay_93_fullRound;
    io_input_payload_delay_94_partialRound <= io_input_payload_delay_93_partialRound;
    io_input_payload_delay_94_stateIndex <= io_input_payload_delay_93_stateIndex;
    io_input_payload_delay_94_stateSize <= io_input_payload_delay_93_stateSize;
    io_input_payload_delay_94_stateID <= io_input_payload_delay_93_stateID;
    io_input_payload_delay_94_stateElements_0 <= io_input_payload_delay_93_stateElements_0;
    io_input_payload_delay_94_stateElements_1 <= io_input_payload_delay_93_stateElements_1;
    io_input_payload_delay_94_stateElements_2 <= io_input_payload_delay_93_stateElements_2;
    io_input_payload_delay_94_stateElements_3 <= io_input_payload_delay_93_stateElements_3;
    io_input_payload_delay_94_stateElements_4 <= io_input_payload_delay_93_stateElements_4;
    io_input_payload_delay_94_stateElements_5 <= io_input_payload_delay_93_stateElements_5;
    io_input_payload_delay_94_stateElements_6 <= io_input_payload_delay_93_stateElements_6;
    io_input_payload_delay_94_stateElements_7 <= io_input_payload_delay_93_stateElements_7;
    io_input_payload_delay_94_stateElements_8 <= io_input_payload_delay_93_stateElements_8;
    io_input_payload_delay_94_stateElements_9 <= io_input_payload_delay_93_stateElements_9;
    io_input_payload_delay_94_stateElements_10 <= io_input_payload_delay_93_stateElements_10;
    io_input_payload_delay_94_stateElement <= io_input_payload_delay_93_stateElement;
    io_input_payload_delay_95_isFull <= io_input_payload_delay_94_isFull;
    io_input_payload_delay_95_fullRound <= io_input_payload_delay_94_fullRound;
    io_input_payload_delay_95_partialRound <= io_input_payload_delay_94_partialRound;
    io_input_payload_delay_95_stateIndex <= io_input_payload_delay_94_stateIndex;
    io_input_payload_delay_95_stateSize <= io_input_payload_delay_94_stateSize;
    io_input_payload_delay_95_stateID <= io_input_payload_delay_94_stateID;
    io_input_payload_delay_95_stateElements_0 <= io_input_payload_delay_94_stateElements_0;
    io_input_payload_delay_95_stateElements_1 <= io_input_payload_delay_94_stateElements_1;
    io_input_payload_delay_95_stateElements_2 <= io_input_payload_delay_94_stateElements_2;
    io_input_payload_delay_95_stateElements_3 <= io_input_payload_delay_94_stateElements_3;
    io_input_payload_delay_95_stateElements_4 <= io_input_payload_delay_94_stateElements_4;
    io_input_payload_delay_95_stateElements_5 <= io_input_payload_delay_94_stateElements_5;
    io_input_payload_delay_95_stateElements_6 <= io_input_payload_delay_94_stateElements_6;
    io_input_payload_delay_95_stateElements_7 <= io_input_payload_delay_94_stateElements_7;
    io_input_payload_delay_95_stateElements_8 <= io_input_payload_delay_94_stateElements_8;
    io_input_payload_delay_95_stateElements_9 <= io_input_payload_delay_94_stateElements_9;
    io_input_payload_delay_95_stateElements_10 <= io_input_payload_delay_94_stateElements_10;
    io_input_payload_delay_95_stateElement <= io_input_payload_delay_94_stateElement;
    io_input_payload_delay_96_isFull <= io_input_payload_delay_95_isFull;
    io_input_payload_delay_96_fullRound <= io_input_payload_delay_95_fullRound;
    io_input_payload_delay_96_partialRound <= io_input_payload_delay_95_partialRound;
    io_input_payload_delay_96_stateIndex <= io_input_payload_delay_95_stateIndex;
    io_input_payload_delay_96_stateSize <= io_input_payload_delay_95_stateSize;
    io_input_payload_delay_96_stateID <= io_input_payload_delay_95_stateID;
    io_input_payload_delay_96_stateElements_0 <= io_input_payload_delay_95_stateElements_0;
    io_input_payload_delay_96_stateElements_1 <= io_input_payload_delay_95_stateElements_1;
    io_input_payload_delay_96_stateElements_2 <= io_input_payload_delay_95_stateElements_2;
    io_input_payload_delay_96_stateElements_3 <= io_input_payload_delay_95_stateElements_3;
    io_input_payload_delay_96_stateElements_4 <= io_input_payload_delay_95_stateElements_4;
    io_input_payload_delay_96_stateElements_5 <= io_input_payload_delay_95_stateElements_5;
    io_input_payload_delay_96_stateElements_6 <= io_input_payload_delay_95_stateElements_6;
    io_input_payload_delay_96_stateElements_7 <= io_input_payload_delay_95_stateElements_7;
    io_input_payload_delay_96_stateElements_8 <= io_input_payload_delay_95_stateElements_8;
    io_input_payload_delay_96_stateElements_9 <= io_input_payload_delay_95_stateElements_9;
    io_input_payload_delay_96_stateElements_10 <= io_input_payload_delay_95_stateElements_10;
    io_input_payload_delay_96_stateElement <= io_input_payload_delay_95_stateElement;
    io_input_payload_delay_97_isFull <= io_input_payload_delay_96_isFull;
    io_input_payload_delay_97_fullRound <= io_input_payload_delay_96_fullRound;
    io_input_payload_delay_97_partialRound <= io_input_payload_delay_96_partialRound;
    io_input_payload_delay_97_stateIndex <= io_input_payload_delay_96_stateIndex;
    io_input_payload_delay_97_stateSize <= io_input_payload_delay_96_stateSize;
    io_input_payload_delay_97_stateID <= io_input_payload_delay_96_stateID;
    io_input_payload_delay_97_stateElements_0 <= io_input_payload_delay_96_stateElements_0;
    io_input_payload_delay_97_stateElements_1 <= io_input_payload_delay_96_stateElements_1;
    io_input_payload_delay_97_stateElements_2 <= io_input_payload_delay_96_stateElements_2;
    io_input_payload_delay_97_stateElements_3 <= io_input_payload_delay_96_stateElements_3;
    io_input_payload_delay_97_stateElements_4 <= io_input_payload_delay_96_stateElements_4;
    io_input_payload_delay_97_stateElements_5 <= io_input_payload_delay_96_stateElements_5;
    io_input_payload_delay_97_stateElements_6 <= io_input_payload_delay_96_stateElements_6;
    io_input_payload_delay_97_stateElements_7 <= io_input_payload_delay_96_stateElements_7;
    io_input_payload_delay_97_stateElements_8 <= io_input_payload_delay_96_stateElements_8;
    io_input_payload_delay_97_stateElements_9 <= io_input_payload_delay_96_stateElements_9;
    io_input_payload_delay_97_stateElements_10 <= io_input_payload_delay_96_stateElements_10;
    io_input_payload_delay_97_stateElement <= io_input_payload_delay_96_stateElement;
    SBox5Stage_tempContext1_isFull <= io_input_payload_delay_97_isFull;
    SBox5Stage_tempContext1_fullRound <= io_input_payload_delay_97_fullRound;
    SBox5Stage_tempContext1_partialRound <= io_input_payload_delay_97_partialRound;
    SBox5Stage_tempContext1_stateIndex <= io_input_payload_delay_97_stateIndex;
    SBox5Stage_tempContext1_stateSize <= io_input_payload_delay_97_stateSize;
    SBox5Stage_tempContext1_stateID <= io_input_payload_delay_97_stateID;
    SBox5Stage_tempContext1_stateElements_0 <= io_input_payload_delay_97_stateElements_0;
    SBox5Stage_tempContext1_stateElements_1 <= io_input_payload_delay_97_stateElements_1;
    SBox5Stage_tempContext1_stateElements_2 <= io_input_payload_delay_97_stateElements_2;
    SBox5Stage_tempContext1_stateElements_3 <= io_input_payload_delay_97_stateElements_3;
    SBox5Stage_tempContext1_stateElements_4 <= io_input_payload_delay_97_stateElements_4;
    SBox5Stage_tempContext1_stateElements_5 <= io_input_payload_delay_97_stateElements_5;
    SBox5Stage_tempContext1_stateElements_6 <= io_input_payload_delay_97_stateElements_6;
    SBox5Stage_tempContext1_stateElements_7 <= io_input_payload_delay_97_stateElements_7;
    SBox5Stage_tempContext1_stateElements_8 <= io_input_payload_delay_97_stateElements_8;
    SBox5Stage_tempContext1_stateElements_9 <= io_input_payload_delay_97_stateElements_9;
    SBox5Stage_tempContext1_stateElements_10 <= io_input_payload_delay_97_stateElements_10;
    SBox5Stage_tempContext1_stateElement <= io_input_payload_delay_97_stateElement;
    SBox5Stage_mul2Context_delay_1_isFull <= SBox5Stage_mul2Context_isFull;
    SBox5Stage_mul2Context_delay_1_fullRound <= SBox5Stage_mul2Context_fullRound;
    SBox5Stage_mul2Context_delay_1_partialRound <= SBox5Stage_mul2Context_partialRound;
    SBox5Stage_mul2Context_delay_1_stateIndex <= SBox5Stage_mul2Context_stateIndex;
    SBox5Stage_mul2Context_delay_1_stateSize <= SBox5Stage_mul2Context_stateSize;
    SBox5Stage_mul2Context_delay_1_stateID <= SBox5Stage_mul2Context_stateID;
    SBox5Stage_mul2Context_delay_1_stateElements_0 <= SBox5Stage_mul2Context_stateElements_0;
    SBox5Stage_mul2Context_delay_1_stateElements_1 <= SBox5Stage_mul2Context_stateElements_1;
    SBox5Stage_mul2Context_delay_1_stateElements_2 <= SBox5Stage_mul2Context_stateElements_2;
    SBox5Stage_mul2Context_delay_1_stateElements_3 <= SBox5Stage_mul2Context_stateElements_3;
    SBox5Stage_mul2Context_delay_1_stateElements_4 <= SBox5Stage_mul2Context_stateElements_4;
    SBox5Stage_mul2Context_delay_1_stateElements_5 <= SBox5Stage_mul2Context_stateElements_5;
    SBox5Stage_mul2Context_delay_1_stateElements_6 <= SBox5Stage_mul2Context_stateElements_6;
    SBox5Stage_mul2Context_delay_1_stateElements_7 <= SBox5Stage_mul2Context_stateElements_7;
    SBox5Stage_mul2Context_delay_1_stateElements_8 <= SBox5Stage_mul2Context_stateElements_8;
    SBox5Stage_mul2Context_delay_1_stateElements_9 <= SBox5Stage_mul2Context_stateElements_9;
    SBox5Stage_mul2Context_delay_1_stateElements_10 <= SBox5Stage_mul2Context_stateElements_10;
    SBox5Stage_mul2Context_delay_2_isFull <= SBox5Stage_mul2Context_delay_1_isFull;
    SBox5Stage_mul2Context_delay_2_fullRound <= SBox5Stage_mul2Context_delay_1_fullRound;
    SBox5Stage_mul2Context_delay_2_partialRound <= SBox5Stage_mul2Context_delay_1_partialRound;
    SBox5Stage_mul2Context_delay_2_stateIndex <= SBox5Stage_mul2Context_delay_1_stateIndex;
    SBox5Stage_mul2Context_delay_2_stateSize <= SBox5Stage_mul2Context_delay_1_stateSize;
    SBox5Stage_mul2Context_delay_2_stateID <= SBox5Stage_mul2Context_delay_1_stateID;
    SBox5Stage_mul2Context_delay_2_stateElements_0 <= SBox5Stage_mul2Context_delay_1_stateElements_0;
    SBox5Stage_mul2Context_delay_2_stateElements_1 <= SBox5Stage_mul2Context_delay_1_stateElements_1;
    SBox5Stage_mul2Context_delay_2_stateElements_2 <= SBox5Stage_mul2Context_delay_1_stateElements_2;
    SBox5Stage_mul2Context_delay_2_stateElements_3 <= SBox5Stage_mul2Context_delay_1_stateElements_3;
    SBox5Stage_mul2Context_delay_2_stateElements_4 <= SBox5Stage_mul2Context_delay_1_stateElements_4;
    SBox5Stage_mul2Context_delay_2_stateElements_5 <= SBox5Stage_mul2Context_delay_1_stateElements_5;
    SBox5Stage_mul2Context_delay_2_stateElements_6 <= SBox5Stage_mul2Context_delay_1_stateElements_6;
    SBox5Stage_mul2Context_delay_2_stateElements_7 <= SBox5Stage_mul2Context_delay_1_stateElements_7;
    SBox5Stage_mul2Context_delay_2_stateElements_8 <= SBox5Stage_mul2Context_delay_1_stateElements_8;
    SBox5Stage_mul2Context_delay_2_stateElements_9 <= SBox5Stage_mul2Context_delay_1_stateElements_9;
    SBox5Stage_mul2Context_delay_2_stateElements_10 <= SBox5Stage_mul2Context_delay_1_stateElements_10;
    SBox5Stage_mul2Context_delay_3_isFull <= SBox5Stage_mul2Context_delay_2_isFull;
    SBox5Stage_mul2Context_delay_3_fullRound <= SBox5Stage_mul2Context_delay_2_fullRound;
    SBox5Stage_mul2Context_delay_3_partialRound <= SBox5Stage_mul2Context_delay_2_partialRound;
    SBox5Stage_mul2Context_delay_3_stateIndex <= SBox5Stage_mul2Context_delay_2_stateIndex;
    SBox5Stage_mul2Context_delay_3_stateSize <= SBox5Stage_mul2Context_delay_2_stateSize;
    SBox5Stage_mul2Context_delay_3_stateID <= SBox5Stage_mul2Context_delay_2_stateID;
    SBox5Stage_mul2Context_delay_3_stateElements_0 <= SBox5Stage_mul2Context_delay_2_stateElements_0;
    SBox5Stage_mul2Context_delay_3_stateElements_1 <= SBox5Stage_mul2Context_delay_2_stateElements_1;
    SBox5Stage_mul2Context_delay_3_stateElements_2 <= SBox5Stage_mul2Context_delay_2_stateElements_2;
    SBox5Stage_mul2Context_delay_3_stateElements_3 <= SBox5Stage_mul2Context_delay_2_stateElements_3;
    SBox5Stage_mul2Context_delay_3_stateElements_4 <= SBox5Stage_mul2Context_delay_2_stateElements_4;
    SBox5Stage_mul2Context_delay_3_stateElements_5 <= SBox5Stage_mul2Context_delay_2_stateElements_5;
    SBox5Stage_mul2Context_delay_3_stateElements_6 <= SBox5Stage_mul2Context_delay_2_stateElements_6;
    SBox5Stage_mul2Context_delay_3_stateElements_7 <= SBox5Stage_mul2Context_delay_2_stateElements_7;
    SBox5Stage_mul2Context_delay_3_stateElements_8 <= SBox5Stage_mul2Context_delay_2_stateElements_8;
    SBox5Stage_mul2Context_delay_3_stateElements_9 <= SBox5Stage_mul2Context_delay_2_stateElements_9;
    SBox5Stage_mul2Context_delay_3_stateElements_10 <= SBox5Stage_mul2Context_delay_2_stateElements_10;
    SBox5Stage_mul2Context_delay_4_isFull <= SBox5Stage_mul2Context_delay_3_isFull;
    SBox5Stage_mul2Context_delay_4_fullRound <= SBox5Stage_mul2Context_delay_3_fullRound;
    SBox5Stage_mul2Context_delay_4_partialRound <= SBox5Stage_mul2Context_delay_3_partialRound;
    SBox5Stage_mul2Context_delay_4_stateIndex <= SBox5Stage_mul2Context_delay_3_stateIndex;
    SBox5Stage_mul2Context_delay_4_stateSize <= SBox5Stage_mul2Context_delay_3_stateSize;
    SBox5Stage_mul2Context_delay_4_stateID <= SBox5Stage_mul2Context_delay_3_stateID;
    SBox5Stage_mul2Context_delay_4_stateElements_0 <= SBox5Stage_mul2Context_delay_3_stateElements_0;
    SBox5Stage_mul2Context_delay_4_stateElements_1 <= SBox5Stage_mul2Context_delay_3_stateElements_1;
    SBox5Stage_mul2Context_delay_4_stateElements_2 <= SBox5Stage_mul2Context_delay_3_stateElements_2;
    SBox5Stage_mul2Context_delay_4_stateElements_3 <= SBox5Stage_mul2Context_delay_3_stateElements_3;
    SBox5Stage_mul2Context_delay_4_stateElements_4 <= SBox5Stage_mul2Context_delay_3_stateElements_4;
    SBox5Stage_mul2Context_delay_4_stateElements_5 <= SBox5Stage_mul2Context_delay_3_stateElements_5;
    SBox5Stage_mul2Context_delay_4_stateElements_6 <= SBox5Stage_mul2Context_delay_3_stateElements_6;
    SBox5Stage_mul2Context_delay_4_stateElements_7 <= SBox5Stage_mul2Context_delay_3_stateElements_7;
    SBox5Stage_mul2Context_delay_4_stateElements_8 <= SBox5Stage_mul2Context_delay_3_stateElements_8;
    SBox5Stage_mul2Context_delay_4_stateElements_9 <= SBox5Stage_mul2Context_delay_3_stateElements_9;
    SBox5Stage_mul2Context_delay_4_stateElements_10 <= SBox5Stage_mul2Context_delay_3_stateElements_10;
    SBox5Stage_mul2Context_delay_5_isFull <= SBox5Stage_mul2Context_delay_4_isFull;
    SBox5Stage_mul2Context_delay_5_fullRound <= SBox5Stage_mul2Context_delay_4_fullRound;
    SBox5Stage_mul2Context_delay_5_partialRound <= SBox5Stage_mul2Context_delay_4_partialRound;
    SBox5Stage_mul2Context_delay_5_stateIndex <= SBox5Stage_mul2Context_delay_4_stateIndex;
    SBox5Stage_mul2Context_delay_5_stateSize <= SBox5Stage_mul2Context_delay_4_stateSize;
    SBox5Stage_mul2Context_delay_5_stateID <= SBox5Stage_mul2Context_delay_4_stateID;
    SBox5Stage_mul2Context_delay_5_stateElements_0 <= SBox5Stage_mul2Context_delay_4_stateElements_0;
    SBox5Stage_mul2Context_delay_5_stateElements_1 <= SBox5Stage_mul2Context_delay_4_stateElements_1;
    SBox5Stage_mul2Context_delay_5_stateElements_2 <= SBox5Stage_mul2Context_delay_4_stateElements_2;
    SBox5Stage_mul2Context_delay_5_stateElements_3 <= SBox5Stage_mul2Context_delay_4_stateElements_3;
    SBox5Stage_mul2Context_delay_5_stateElements_4 <= SBox5Stage_mul2Context_delay_4_stateElements_4;
    SBox5Stage_mul2Context_delay_5_stateElements_5 <= SBox5Stage_mul2Context_delay_4_stateElements_5;
    SBox5Stage_mul2Context_delay_5_stateElements_6 <= SBox5Stage_mul2Context_delay_4_stateElements_6;
    SBox5Stage_mul2Context_delay_5_stateElements_7 <= SBox5Stage_mul2Context_delay_4_stateElements_7;
    SBox5Stage_mul2Context_delay_5_stateElements_8 <= SBox5Stage_mul2Context_delay_4_stateElements_8;
    SBox5Stage_mul2Context_delay_5_stateElements_9 <= SBox5Stage_mul2Context_delay_4_stateElements_9;
    SBox5Stage_mul2Context_delay_5_stateElements_10 <= SBox5Stage_mul2Context_delay_4_stateElements_10;
    SBox5Stage_mul2Context_delay_6_isFull <= SBox5Stage_mul2Context_delay_5_isFull;
    SBox5Stage_mul2Context_delay_6_fullRound <= SBox5Stage_mul2Context_delay_5_fullRound;
    SBox5Stage_mul2Context_delay_6_partialRound <= SBox5Stage_mul2Context_delay_5_partialRound;
    SBox5Stage_mul2Context_delay_6_stateIndex <= SBox5Stage_mul2Context_delay_5_stateIndex;
    SBox5Stage_mul2Context_delay_6_stateSize <= SBox5Stage_mul2Context_delay_5_stateSize;
    SBox5Stage_mul2Context_delay_6_stateID <= SBox5Stage_mul2Context_delay_5_stateID;
    SBox5Stage_mul2Context_delay_6_stateElements_0 <= SBox5Stage_mul2Context_delay_5_stateElements_0;
    SBox5Stage_mul2Context_delay_6_stateElements_1 <= SBox5Stage_mul2Context_delay_5_stateElements_1;
    SBox5Stage_mul2Context_delay_6_stateElements_2 <= SBox5Stage_mul2Context_delay_5_stateElements_2;
    SBox5Stage_mul2Context_delay_6_stateElements_3 <= SBox5Stage_mul2Context_delay_5_stateElements_3;
    SBox5Stage_mul2Context_delay_6_stateElements_4 <= SBox5Stage_mul2Context_delay_5_stateElements_4;
    SBox5Stage_mul2Context_delay_6_stateElements_5 <= SBox5Stage_mul2Context_delay_5_stateElements_5;
    SBox5Stage_mul2Context_delay_6_stateElements_6 <= SBox5Stage_mul2Context_delay_5_stateElements_6;
    SBox5Stage_mul2Context_delay_6_stateElements_7 <= SBox5Stage_mul2Context_delay_5_stateElements_7;
    SBox5Stage_mul2Context_delay_6_stateElements_8 <= SBox5Stage_mul2Context_delay_5_stateElements_8;
    SBox5Stage_mul2Context_delay_6_stateElements_9 <= SBox5Stage_mul2Context_delay_5_stateElements_9;
    SBox5Stage_mul2Context_delay_6_stateElements_10 <= SBox5Stage_mul2Context_delay_5_stateElements_10;
    SBox5Stage_mul2Context_delay_7_isFull <= SBox5Stage_mul2Context_delay_6_isFull;
    SBox5Stage_mul2Context_delay_7_fullRound <= SBox5Stage_mul2Context_delay_6_fullRound;
    SBox5Stage_mul2Context_delay_7_partialRound <= SBox5Stage_mul2Context_delay_6_partialRound;
    SBox5Stage_mul2Context_delay_7_stateIndex <= SBox5Stage_mul2Context_delay_6_stateIndex;
    SBox5Stage_mul2Context_delay_7_stateSize <= SBox5Stage_mul2Context_delay_6_stateSize;
    SBox5Stage_mul2Context_delay_7_stateID <= SBox5Stage_mul2Context_delay_6_stateID;
    SBox5Stage_mul2Context_delay_7_stateElements_0 <= SBox5Stage_mul2Context_delay_6_stateElements_0;
    SBox5Stage_mul2Context_delay_7_stateElements_1 <= SBox5Stage_mul2Context_delay_6_stateElements_1;
    SBox5Stage_mul2Context_delay_7_stateElements_2 <= SBox5Stage_mul2Context_delay_6_stateElements_2;
    SBox5Stage_mul2Context_delay_7_stateElements_3 <= SBox5Stage_mul2Context_delay_6_stateElements_3;
    SBox5Stage_mul2Context_delay_7_stateElements_4 <= SBox5Stage_mul2Context_delay_6_stateElements_4;
    SBox5Stage_mul2Context_delay_7_stateElements_5 <= SBox5Stage_mul2Context_delay_6_stateElements_5;
    SBox5Stage_mul2Context_delay_7_stateElements_6 <= SBox5Stage_mul2Context_delay_6_stateElements_6;
    SBox5Stage_mul2Context_delay_7_stateElements_7 <= SBox5Stage_mul2Context_delay_6_stateElements_7;
    SBox5Stage_mul2Context_delay_7_stateElements_8 <= SBox5Stage_mul2Context_delay_6_stateElements_8;
    SBox5Stage_mul2Context_delay_7_stateElements_9 <= SBox5Stage_mul2Context_delay_6_stateElements_9;
    SBox5Stage_mul2Context_delay_7_stateElements_10 <= SBox5Stage_mul2Context_delay_6_stateElements_10;
    SBox5Stage_mul2Context_delay_8_isFull <= SBox5Stage_mul2Context_delay_7_isFull;
    SBox5Stage_mul2Context_delay_8_fullRound <= SBox5Stage_mul2Context_delay_7_fullRound;
    SBox5Stage_mul2Context_delay_8_partialRound <= SBox5Stage_mul2Context_delay_7_partialRound;
    SBox5Stage_mul2Context_delay_8_stateIndex <= SBox5Stage_mul2Context_delay_7_stateIndex;
    SBox5Stage_mul2Context_delay_8_stateSize <= SBox5Stage_mul2Context_delay_7_stateSize;
    SBox5Stage_mul2Context_delay_8_stateID <= SBox5Stage_mul2Context_delay_7_stateID;
    SBox5Stage_mul2Context_delay_8_stateElements_0 <= SBox5Stage_mul2Context_delay_7_stateElements_0;
    SBox5Stage_mul2Context_delay_8_stateElements_1 <= SBox5Stage_mul2Context_delay_7_stateElements_1;
    SBox5Stage_mul2Context_delay_8_stateElements_2 <= SBox5Stage_mul2Context_delay_7_stateElements_2;
    SBox5Stage_mul2Context_delay_8_stateElements_3 <= SBox5Stage_mul2Context_delay_7_stateElements_3;
    SBox5Stage_mul2Context_delay_8_stateElements_4 <= SBox5Stage_mul2Context_delay_7_stateElements_4;
    SBox5Stage_mul2Context_delay_8_stateElements_5 <= SBox5Stage_mul2Context_delay_7_stateElements_5;
    SBox5Stage_mul2Context_delay_8_stateElements_6 <= SBox5Stage_mul2Context_delay_7_stateElements_6;
    SBox5Stage_mul2Context_delay_8_stateElements_7 <= SBox5Stage_mul2Context_delay_7_stateElements_7;
    SBox5Stage_mul2Context_delay_8_stateElements_8 <= SBox5Stage_mul2Context_delay_7_stateElements_8;
    SBox5Stage_mul2Context_delay_8_stateElements_9 <= SBox5Stage_mul2Context_delay_7_stateElements_9;
    SBox5Stage_mul2Context_delay_8_stateElements_10 <= SBox5Stage_mul2Context_delay_7_stateElements_10;
    SBox5Stage_mul2Context_delay_9_isFull <= SBox5Stage_mul2Context_delay_8_isFull;
    SBox5Stage_mul2Context_delay_9_fullRound <= SBox5Stage_mul2Context_delay_8_fullRound;
    SBox5Stage_mul2Context_delay_9_partialRound <= SBox5Stage_mul2Context_delay_8_partialRound;
    SBox5Stage_mul2Context_delay_9_stateIndex <= SBox5Stage_mul2Context_delay_8_stateIndex;
    SBox5Stage_mul2Context_delay_9_stateSize <= SBox5Stage_mul2Context_delay_8_stateSize;
    SBox5Stage_mul2Context_delay_9_stateID <= SBox5Stage_mul2Context_delay_8_stateID;
    SBox5Stage_mul2Context_delay_9_stateElements_0 <= SBox5Stage_mul2Context_delay_8_stateElements_0;
    SBox5Stage_mul2Context_delay_9_stateElements_1 <= SBox5Stage_mul2Context_delay_8_stateElements_1;
    SBox5Stage_mul2Context_delay_9_stateElements_2 <= SBox5Stage_mul2Context_delay_8_stateElements_2;
    SBox5Stage_mul2Context_delay_9_stateElements_3 <= SBox5Stage_mul2Context_delay_8_stateElements_3;
    SBox5Stage_mul2Context_delay_9_stateElements_4 <= SBox5Stage_mul2Context_delay_8_stateElements_4;
    SBox5Stage_mul2Context_delay_9_stateElements_5 <= SBox5Stage_mul2Context_delay_8_stateElements_5;
    SBox5Stage_mul2Context_delay_9_stateElements_6 <= SBox5Stage_mul2Context_delay_8_stateElements_6;
    SBox5Stage_mul2Context_delay_9_stateElements_7 <= SBox5Stage_mul2Context_delay_8_stateElements_7;
    SBox5Stage_mul2Context_delay_9_stateElements_8 <= SBox5Stage_mul2Context_delay_8_stateElements_8;
    SBox5Stage_mul2Context_delay_9_stateElements_9 <= SBox5Stage_mul2Context_delay_8_stateElements_9;
    SBox5Stage_mul2Context_delay_9_stateElements_10 <= SBox5Stage_mul2Context_delay_8_stateElements_10;
    SBox5Stage_mul2Context_delay_10_isFull <= SBox5Stage_mul2Context_delay_9_isFull;
    SBox5Stage_mul2Context_delay_10_fullRound <= SBox5Stage_mul2Context_delay_9_fullRound;
    SBox5Stage_mul2Context_delay_10_partialRound <= SBox5Stage_mul2Context_delay_9_partialRound;
    SBox5Stage_mul2Context_delay_10_stateIndex <= SBox5Stage_mul2Context_delay_9_stateIndex;
    SBox5Stage_mul2Context_delay_10_stateSize <= SBox5Stage_mul2Context_delay_9_stateSize;
    SBox5Stage_mul2Context_delay_10_stateID <= SBox5Stage_mul2Context_delay_9_stateID;
    SBox5Stage_mul2Context_delay_10_stateElements_0 <= SBox5Stage_mul2Context_delay_9_stateElements_0;
    SBox5Stage_mul2Context_delay_10_stateElements_1 <= SBox5Stage_mul2Context_delay_9_stateElements_1;
    SBox5Stage_mul2Context_delay_10_stateElements_2 <= SBox5Stage_mul2Context_delay_9_stateElements_2;
    SBox5Stage_mul2Context_delay_10_stateElements_3 <= SBox5Stage_mul2Context_delay_9_stateElements_3;
    SBox5Stage_mul2Context_delay_10_stateElements_4 <= SBox5Stage_mul2Context_delay_9_stateElements_4;
    SBox5Stage_mul2Context_delay_10_stateElements_5 <= SBox5Stage_mul2Context_delay_9_stateElements_5;
    SBox5Stage_mul2Context_delay_10_stateElements_6 <= SBox5Stage_mul2Context_delay_9_stateElements_6;
    SBox5Stage_mul2Context_delay_10_stateElements_7 <= SBox5Stage_mul2Context_delay_9_stateElements_7;
    SBox5Stage_mul2Context_delay_10_stateElements_8 <= SBox5Stage_mul2Context_delay_9_stateElements_8;
    SBox5Stage_mul2Context_delay_10_stateElements_9 <= SBox5Stage_mul2Context_delay_9_stateElements_9;
    SBox5Stage_mul2Context_delay_10_stateElements_10 <= SBox5Stage_mul2Context_delay_9_stateElements_10;
    SBox5Stage_mul2Context_delay_11_isFull <= SBox5Stage_mul2Context_delay_10_isFull;
    SBox5Stage_mul2Context_delay_11_fullRound <= SBox5Stage_mul2Context_delay_10_fullRound;
    SBox5Stage_mul2Context_delay_11_partialRound <= SBox5Stage_mul2Context_delay_10_partialRound;
    SBox5Stage_mul2Context_delay_11_stateIndex <= SBox5Stage_mul2Context_delay_10_stateIndex;
    SBox5Stage_mul2Context_delay_11_stateSize <= SBox5Stage_mul2Context_delay_10_stateSize;
    SBox5Stage_mul2Context_delay_11_stateID <= SBox5Stage_mul2Context_delay_10_stateID;
    SBox5Stage_mul2Context_delay_11_stateElements_0 <= SBox5Stage_mul2Context_delay_10_stateElements_0;
    SBox5Stage_mul2Context_delay_11_stateElements_1 <= SBox5Stage_mul2Context_delay_10_stateElements_1;
    SBox5Stage_mul2Context_delay_11_stateElements_2 <= SBox5Stage_mul2Context_delay_10_stateElements_2;
    SBox5Stage_mul2Context_delay_11_stateElements_3 <= SBox5Stage_mul2Context_delay_10_stateElements_3;
    SBox5Stage_mul2Context_delay_11_stateElements_4 <= SBox5Stage_mul2Context_delay_10_stateElements_4;
    SBox5Stage_mul2Context_delay_11_stateElements_5 <= SBox5Stage_mul2Context_delay_10_stateElements_5;
    SBox5Stage_mul2Context_delay_11_stateElements_6 <= SBox5Stage_mul2Context_delay_10_stateElements_6;
    SBox5Stage_mul2Context_delay_11_stateElements_7 <= SBox5Stage_mul2Context_delay_10_stateElements_7;
    SBox5Stage_mul2Context_delay_11_stateElements_8 <= SBox5Stage_mul2Context_delay_10_stateElements_8;
    SBox5Stage_mul2Context_delay_11_stateElements_9 <= SBox5Stage_mul2Context_delay_10_stateElements_9;
    SBox5Stage_mul2Context_delay_11_stateElements_10 <= SBox5Stage_mul2Context_delay_10_stateElements_10;
    SBox5Stage_mul2Context_delay_12_isFull <= SBox5Stage_mul2Context_delay_11_isFull;
    SBox5Stage_mul2Context_delay_12_fullRound <= SBox5Stage_mul2Context_delay_11_fullRound;
    SBox5Stage_mul2Context_delay_12_partialRound <= SBox5Stage_mul2Context_delay_11_partialRound;
    SBox5Stage_mul2Context_delay_12_stateIndex <= SBox5Stage_mul2Context_delay_11_stateIndex;
    SBox5Stage_mul2Context_delay_12_stateSize <= SBox5Stage_mul2Context_delay_11_stateSize;
    SBox5Stage_mul2Context_delay_12_stateID <= SBox5Stage_mul2Context_delay_11_stateID;
    SBox5Stage_mul2Context_delay_12_stateElements_0 <= SBox5Stage_mul2Context_delay_11_stateElements_0;
    SBox5Stage_mul2Context_delay_12_stateElements_1 <= SBox5Stage_mul2Context_delay_11_stateElements_1;
    SBox5Stage_mul2Context_delay_12_stateElements_2 <= SBox5Stage_mul2Context_delay_11_stateElements_2;
    SBox5Stage_mul2Context_delay_12_stateElements_3 <= SBox5Stage_mul2Context_delay_11_stateElements_3;
    SBox5Stage_mul2Context_delay_12_stateElements_4 <= SBox5Stage_mul2Context_delay_11_stateElements_4;
    SBox5Stage_mul2Context_delay_12_stateElements_5 <= SBox5Stage_mul2Context_delay_11_stateElements_5;
    SBox5Stage_mul2Context_delay_12_stateElements_6 <= SBox5Stage_mul2Context_delay_11_stateElements_6;
    SBox5Stage_mul2Context_delay_12_stateElements_7 <= SBox5Stage_mul2Context_delay_11_stateElements_7;
    SBox5Stage_mul2Context_delay_12_stateElements_8 <= SBox5Stage_mul2Context_delay_11_stateElements_8;
    SBox5Stage_mul2Context_delay_12_stateElements_9 <= SBox5Stage_mul2Context_delay_11_stateElements_9;
    SBox5Stage_mul2Context_delay_12_stateElements_10 <= SBox5Stage_mul2Context_delay_11_stateElements_10;
    SBox5Stage_mul2Context_delay_13_isFull <= SBox5Stage_mul2Context_delay_12_isFull;
    SBox5Stage_mul2Context_delay_13_fullRound <= SBox5Stage_mul2Context_delay_12_fullRound;
    SBox5Stage_mul2Context_delay_13_partialRound <= SBox5Stage_mul2Context_delay_12_partialRound;
    SBox5Stage_mul2Context_delay_13_stateIndex <= SBox5Stage_mul2Context_delay_12_stateIndex;
    SBox5Stage_mul2Context_delay_13_stateSize <= SBox5Stage_mul2Context_delay_12_stateSize;
    SBox5Stage_mul2Context_delay_13_stateID <= SBox5Stage_mul2Context_delay_12_stateID;
    SBox5Stage_mul2Context_delay_13_stateElements_0 <= SBox5Stage_mul2Context_delay_12_stateElements_0;
    SBox5Stage_mul2Context_delay_13_stateElements_1 <= SBox5Stage_mul2Context_delay_12_stateElements_1;
    SBox5Stage_mul2Context_delay_13_stateElements_2 <= SBox5Stage_mul2Context_delay_12_stateElements_2;
    SBox5Stage_mul2Context_delay_13_stateElements_3 <= SBox5Stage_mul2Context_delay_12_stateElements_3;
    SBox5Stage_mul2Context_delay_13_stateElements_4 <= SBox5Stage_mul2Context_delay_12_stateElements_4;
    SBox5Stage_mul2Context_delay_13_stateElements_5 <= SBox5Stage_mul2Context_delay_12_stateElements_5;
    SBox5Stage_mul2Context_delay_13_stateElements_6 <= SBox5Stage_mul2Context_delay_12_stateElements_6;
    SBox5Stage_mul2Context_delay_13_stateElements_7 <= SBox5Stage_mul2Context_delay_12_stateElements_7;
    SBox5Stage_mul2Context_delay_13_stateElements_8 <= SBox5Stage_mul2Context_delay_12_stateElements_8;
    SBox5Stage_mul2Context_delay_13_stateElements_9 <= SBox5Stage_mul2Context_delay_12_stateElements_9;
    SBox5Stage_mul2Context_delay_13_stateElements_10 <= SBox5Stage_mul2Context_delay_12_stateElements_10;
    SBox5Stage_mul2Context_delay_14_isFull <= SBox5Stage_mul2Context_delay_13_isFull;
    SBox5Stage_mul2Context_delay_14_fullRound <= SBox5Stage_mul2Context_delay_13_fullRound;
    SBox5Stage_mul2Context_delay_14_partialRound <= SBox5Stage_mul2Context_delay_13_partialRound;
    SBox5Stage_mul2Context_delay_14_stateIndex <= SBox5Stage_mul2Context_delay_13_stateIndex;
    SBox5Stage_mul2Context_delay_14_stateSize <= SBox5Stage_mul2Context_delay_13_stateSize;
    SBox5Stage_mul2Context_delay_14_stateID <= SBox5Stage_mul2Context_delay_13_stateID;
    SBox5Stage_mul2Context_delay_14_stateElements_0 <= SBox5Stage_mul2Context_delay_13_stateElements_0;
    SBox5Stage_mul2Context_delay_14_stateElements_1 <= SBox5Stage_mul2Context_delay_13_stateElements_1;
    SBox5Stage_mul2Context_delay_14_stateElements_2 <= SBox5Stage_mul2Context_delay_13_stateElements_2;
    SBox5Stage_mul2Context_delay_14_stateElements_3 <= SBox5Stage_mul2Context_delay_13_stateElements_3;
    SBox5Stage_mul2Context_delay_14_stateElements_4 <= SBox5Stage_mul2Context_delay_13_stateElements_4;
    SBox5Stage_mul2Context_delay_14_stateElements_5 <= SBox5Stage_mul2Context_delay_13_stateElements_5;
    SBox5Stage_mul2Context_delay_14_stateElements_6 <= SBox5Stage_mul2Context_delay_13_stateElements_6;
    SBox5Stage_mul2Context_delay_14_stateElements_7 <= SBox5Stage_mul2Context_delay_13_stateElements_7;
    SBox5Stage_mul2Context_delay_14_stateElements_8 <= SBox5Stage_mul2Context_delay_13_stateElements_8;
    SBox5Stage_mul2Context_delay_14_stateElements_9 <= SBox5Stage_mul2Context_delay_13_stateElements_9;
    SBox5Stage_mul2Context_delay_14_stateElements_10 <= SBox5Stage_mul2Context_delay_13_stateElements_10;
    SBox5Stage_mul2Context_delay_15_isFull <= SBox5Stage_mul2Context_delay_14_isFull;
    SBox5Stage_mul2Context_delay_15_fullRound <= SBox5Stage_mul2Context_delay_14_fullRound;
    SBox5Stage_mul2Context_delay_15_partialRound <= SBox5Stage_mul2Context_delay_14_partialRound;
    SBox5Stage_mul2Context_delay_15_stateIndex <= SBox5Stage_mul2Context_delay_14_stateIndex;
    SBox5Stage_mul2Context_delay_15_stateSize <= SBox5Stage_mul2Context_delay_14_stateSize;
    SBox5Stage_mul2Context_delay_15_stateID <= SBox5Stage_mul2Context_delay_14_stateID;
    SBox5Stage_mul2Context_delay_15_stateElements_0 <= SBox5Stage_mul2Context_delay_14_stateElements_0;
    SBox5Stage_mul2Context_delay_15_stateElements_1 <= SBox5Stage_mul2Context_delay_14_stateElements_1;
    SBox5Stage_mul2Context_delay_15_stateElements_2 <= SBox5Stage_mul2Context_delay_14_stateElements_2;
    SBox5Stage_mul2Context_delay_15_stateElements_3 <= SBox5Stage_mul2Context_delay_14_stateElements_3;
    SBox5Stage_mul2Context_delay_15_stateElements_4 <= SBox5Stage_mul2Context_delay_14_stateElements_4;
    SBox5Stage_mul2Context_delay_15_stateElements_5 <= SBox5Stage_mul2Context_delay_14_stateElements_5;
    SBox5Stage_mul2Context_delay_15_stateElements_6 <= SBox5Stage_mul2Context_delay_14_stateElements_6;
    SBox5Stage_mul2Context_delay_15_stateElements_7 <= SBox5Stage_mul2Context_delay_14_stateElements_7;
    SBox5Stage_mul2Context_delay_15_stateElements_8 <= SBox5Stage_mul2Context_delay_14_stateElements_8;
    SBox5Stage_mul2Context_delay_15_stateElements_9 <= SBox5Stage_mul2Context_delay_14_stateElements_9;
    SBox5Stage_mul2Context_delay_15_stateElements_10 <= SBox5Stage_mul2Context_delay_14_stateElements_10;
    SBox5Stage_mul2Context_delay_16_isFull <= SBox5Stage_mul2Context_delay_15_isFull;
    SBox5Stage_mul2Context_delay_16_fullRound <= SBox5Stage_mul2Context_delay_15_fullRound;
    SBox5Stage_mul2Context_delay_16_partialRound <= SBox5Stage_mul2Context_delay_15_partialRound;
    SBox5Stage_mul2Context_delay_16_stateIndex <= SBox5Stage_mul2Context_delay_15_stateIndex;
    SBox5Stage_mul2Context_delay_16_stateSize <= SBox5Stage_mul2Context_delay_15_stateSize;
    SBox5Stage_mul2Context_delay_16_stateID <= SBox5Stage_mul2Context_delay_15_stateID;
    SBox5Stage_mul2Context_delay_16_stateElements_0 <= SBox5Stage_mul2Context_delay_15_stateElements_0;
    SBox5Stage_mul2Context_delay_16_stateElements_1 <= SBox5Stage_mul2Context_delay_15_stateElements_1;
    SBox5Stage_mul2Context_delay_16_stateElements_2 <= SBox5Stage_mul2Context_delay_15_stateElements_2;
    SBox5Stage_mul2Context_delay_16_stateElements_3 <= SBox5Stage_mul2Context_delay_15_stateElements_3;
    SBox5Stage_mul2Context_delay_16_stateElements_4 <= SBox5Stage_mul2Context_delay_15_stateElements_4;
    SBox5Stage_mul2Context_delay_16_stateElements_5 <= SBox5Stage_mul2Context_delay_15_stateElements_5;
    SBox5Stage_mul2Context_delay_16_stateElements_6 <= SBox5Stage_mul2Context_delay_15_stateElements_6;
    SBox5Stage_mul2Context_delay_16_stateElements_7 <= SBox5Stage_mul2Context_delay_15_stateElements_7;
    SBox5Stage_mul2Context_delay_16_stateElements_8 <= SBox5Stage_mul2Context_delay_15_stateElements_8;
    SBox5Stage_mul2Context_delay_16_stateElements_9 <= SBox5Stage_mul2Context_delay_15_stateElements_9;
    SBox5Stage_mul2Context_delay_16_stateElements_10 <= SBox5Stage_mul2Context_delay_15_stateElements_10;
    SBox5Stage_mul2Context_delay_17_isFull <= SBox5Stage_mul2Context_delay_16_isFull;
    SBox5Stage_mul2Context_delay_17_fullRound <= SBox5Stage_mul2Context_delay_16_fullRound;
    SBox5Stage_mul2Context_delay_17_partialRound <= SBox5Stage_mul2Context_delay_16_partialRound;
    SBox5Stage_mul2Context_delay_17_stateIndex <= SBox5Stage_mul2Context_delay_16_stateIndex;
    SBox5Stage_mul2Context_delay_17_stateSize <= SBox5Stage_mul2Context_delay_16_stateSize;
    SBox5Stage_mul2Context_delay_17_stateID <= SBox5Stage_mul2Context_delay_16_stateID;
    SBox5Stage_mul2Context_delay_17_stateElements_0 <= SBox5Stage_mul2Context_delay_16_stateElements_0;
    SBox5Stage_mul2Context_delay_17_stateElements_1 <= SBox5Stage_mul2Context_delay_16_stateElements_1;
    SBox5Stage_mul2Context_delay_17_stateElements_2 <= SBox5Stage_mul2Context_delay_16_stateElements_2;
    SBox5Stage_mul2Context_delay_17_stateElements_3 <= SBox5Stage_mul2Context_delay_16_stateElements_3;
    SBox5Stage_mul2Context_delay_17_stateElements_4 <= SBox5Stage_mul2Context_delay_16_stateElements_4;
    SBox5Stage_mul2Context_delay_17_stateElements_5 <= SBox5Stage_mul2Context_delay_16_stateElements_5;
    SBox5Stage_mul2Context_delay_17_stateElements_6 <= SBox5Stage_mul2Context_delay_16_stateElements_6;
    SBox5Stage_mul2Context_delay_17_stateElements_7 <= SBox5Stage_mul2Context_delay_16_stateElements_7;
    SBox5Stage_mul2Context_delay_17_stateElements_8 <= SBox5Stage_mul2Context_delay_16_stateElements_8;
    SBox5Stage_mul2Context_delay_17_stateElements_9 <= SBox5Stage_mul2Context_delay_16_stateElements_9;
    SBox5Stage_mul2Context_delay_17_stateElements_10 <= SBox5Stage_mul2Context_delay_16_stateElements_10;
    SBox5Stage_mul2Context_delay_18_isFull <= SBox5Stage_mul2Context_delay_17_isFull;
    SBox5Stage_mul2Context_delay_18_fullRound <= SBox5Stage_mul2Context_delay_17_fullRound;
    SBox5Stage_mul2Context_delay_18_partialRound <= SBox5Stage_mul2Context_delay_17_partialRound;
    SBox5Stage_mul2Context_delay_18_stateIndex <= SBox5Stage_mul2Context_delay_17_stateIndex;
    SBox5Stage_mul2Context_delay_18_stateSize <= SBox5Stage_mul2Context_delay_17_stateSize;
    SBox5Stage_mul2Context_delay_18_stateID <= SBox5Stage_mul2Context_delay_17_stateID;
    SBox5Stage_mul2Context_delay_18_stateElements_0 <= SBox5Stage_mul2Context_delay_17_stateElements_0;
    SBox5Stage_mul2Context_delay_18_stateElements_1 <= SBox5Stage_mul2Context_delay_17_stateElements_1;
    SBox5Stage_mul2Context_delay_18_stateElements_2 <= SBox5Stage_mul2Context_delay_17_stateElements_2;
    SBox5Stage_mul2Context_delay_18_stateElements_3 <= SBox5Stage_mul2Context_delay_17_stateElements_3;
    SBox5Stage_mul2Context_delay_18_stateElements_4 <= SBox5Stage_mul2Context_delay_17_stateElements_4;
    SBox5Stage_mul2Context_delay_18_stateElements_5 <= SBox5Stage_mul2Context_delay_17_stateElements_5;
    SBox5Stage_mul2Context_delay_18_stateElements_6 <= SBox5Stage_mul2Context_delay_17_stateElements_6;
    SBox5Stage_mul2Context_delay_18_stateElements_7 <= SBox5Stage_mul2Context_delay_17_stateElements_7;
    SBox5Stage_mul2Context_delay_18_stateElements_8 <= SBox5Stage_mul2Context_delay_17_stateElements_8;
    SBox5Stage_mul2Context_delay_18_stateElements_9 <= SBox5Stage_mul2Context_delay_17_stateElements_9;
    SBox5Stage_mul2Context_delay_18_stateElements_10 <= SBox5Stage_mul2Context_delay_17_stateElements_10;
    SBox5Stage_mul2Context_delay_19_isFull <= SBox5Stage_mul2Context_delay_18_isFull;
    SBox5Stage_mul2Context_delay_19_fullRound <= SBox5Stage_mul2Context_delay_18_fullRound;
    SBox5Stage_mul2Context_delay_19_partialRound <= SBox5Stage_mul2Context_delay_18_partialRound;
    SBox5Stage_mul2Context_delay_19_stateIndex <= SBox5Stage_mul2Context_delay_18_stateIndex;
    SBox5Stage_mul2Context_delay_19_stateSize <= SBox5Stage_mul2Context_delay_18_stateSize;
    SBox5Stage_mul2Context_delay_19_stateID <= SBox5Stage_mul2Context_delay_18_stateID;
    SBox5Stage_mul2Context_delay_19_stateElements_0 <= SBox5Stage_mul2Context_delay_18_stateElements_0;
    SBox5Stage_mul2Context_delay_19_stateElements_1 <= SBox5Stage_mul2Context_delay_18_stateElements_1;
    SBox5Stage_mul2Context_delay_19_stateElements_2 <= SBox5Stage_mul2Context_delay_18_stateElements_2;
    SBox5Stage_mul2Context_delay_19_stateElements_3 <= SBox5Stage_mul2Context_delay_18_stateElements_3;
    SBox5Stage_mul2Context_delay_19_stateElements_4 <= SBox5Stage_mul2Context_delay_18_stateElements_4;
    SBox5Stage_mul2Context_delay_19_stateElements_5 <= SBox5Stage_mul2Context_delay_18_stateElements_5;
    SBox5Stage_mul2Context_delay_19_stateElements_6 <= SBox5Stage_mul2Context_delay_18_stateElements_6;
    SBox5Stage_mul2Context_delay_19_stateElements_7 <= SBox5Stage_mul2Context_delay_18_stateElements_7;
    SBox5Stage_mul2Context_delay_19_stateElements_8 <= SBox5Stage_mul2Context_delay_18_stateElements_8;
    SBox5Stage_mul2Context_delay_19_stateElements_9 <= SBox5Stage_mul2Context_delay_18_stateElements_9;
    SBox5Stage_mul2Context_delay_19_stateElements_10 <= SBox5Stage_mul2Context_delay_18_stateElements_10;
    SBox5Stage_mul2Context_delay_20_isFull <= SBox5Stage_mul2Context_delay_19_isFull;
    SBox5Stage_mul2Context_delay_20_fullRound <= SBox5Stage_mul2Context_delay_19_fullRound;
    SBox5Stage_mul2Context_delay_20_partialRound <= SBox5Stage_mul2Context_delay_19_partialRound;
    SBox5Stage_mul2Context_delay_20_stateIndex <= SBox5Stage_mul2Context_delay_19_stateIndex;
    SBox5Stage_mul2Context_delay_20_stateSize <= SBox5Stage_mul2Context_delay_19_stateSize;
    SBox5Stage_mul2Context_delay_20_stateID <= SBox5Stage_mul2Context_delay_19_stateID;
    SBox5Stage_mul2Context_delay_20_stateElements_0 <= SBox5Stage_mul2Context_delay_19_stateElements_0;
    SBox5Stage_mul2Context_delay_20_stateElements_1 <= SBox5Stage_mul2Context_delay_19_stateElements_1;
    SBox5Stage_mul2Context_delay_20_stateElements_2 <= SBox5Stage_mul2Context_delay_19_stateElements_2;
    SBox5Stage_mul2Context_delay_20_stateElements_3 <= SBox5Stage_mul2Context_delay_19_stateElements_3;
    SBox5Stage_mul2Context_delay_20_stateElements_4 <= SBox5Stage_mul2Context_delay_19_stateElements_4;
    SBox5Stage_mul2Context_delay_20_stateElements_5 <= SBox5Stage_mul2Context_delay_19_stateElements_5;
    SBox5Stage_mul2Context_delay_20_stateElements_6 <= SBox5Stage_mul2Context_delay_19_stateElements_6;
    SBox5Stage_mul2Context_delay_20_stateElements_7 <= SBox5Stage_mul2Context_delay_19_stateElements_7;
    SBox5Stage_mul2Context_delay_20_stateElements_8 <= SBox5Stage_mul2Context_delay_19_stateElements_8;
    SBox5Stage_mul2Context_delay_20_stateElements_9 <= SBox5Stage_mul2Context_delay_19_stateElements_9;
    SBox5Stage_mul2Context_delay_20_stateElements_10 <= SBox5Stage_mul2Context_delay_19_stateElements_10;
    SBox5Stage_mul2Context_delay_21_isFull <= SBox5Stage_mul2Context_delay_20_isFull;
    SBox5Stage_mul2Context_delay_21_fullRound <= SBox5Stage_mul2Context_delay_20_fullRound;
    SBox5Stage_mul2Context_delay_21_partialRound <= SBox5Stage_mul2Context_delay_20_partialRound;
    SBox5Stage_mul2Context_delay_21_stateIndex <= SBox5Stage_mul2Context_delay_20_stateIndex;
    SBox5Stage_mul2Context_delay_21_stateSize <= SBox5Stage_mul2Context_delay_20_stateSize;
    SBox5Stage_mul2Context_delay_21_stateID <= SBox5Stage_mul2Context_delay_20_stateID;
    SBox5Stage_mul2Context_delay_21_stateElements_0 <= SBox5Stage_mul2Context_delay_20_stateElements_0;
    SBox5Stage_mul2Context_delay_21_stateElements_1 <= SBox5Stage_mul2Context_delay_20_stateElements_1;
    SBox5Stage_mul2Context_delay_21_stateElements_2 <= SBox5Stage_mul2Context_delay_20_stateElements_2;
    SBox5Stage_mul2Context_delay_21_stateElements_3 <= SBox5Stage_mul2Context_delay_20_stateElements_3;
    SBox5Stage_mul2Context_delay_21_stateElements_4 <= SBox5Stage_mul2Context_delay_20_stateElements_4;
    SBox5Stage_mul2Context_delay_21_stateElements_5 <= SBox5Stage_mul2Context_delay_20_stateElements_5;
    SBox5Stage_mul2Context_delay_21_stateElements_6 <= SBox5Stage_mul2Context_delay_20_stateElements_6;
    SBox5Stage_mul2Context_delay_21_stateElements_7 <= SBox5Stage_mul2Context_delay_20_stateElements_7;
    SBox5Stage_mul2Context_delay_21_stateElements_8 <= SBox5Stage_mul2Context_delay_20_stateElements_8;
    SBox5Stage_mul2Context_delay_21_stateElements_9 <= SBox5Stage_mul2Context_delay_20_stateElements_9;
    SBox5Stage_mul2Context_delay_21_stateElements_10 <= SBox5Stage_mul2Context_delay_20_stateElements_10;
    SBox5Stage_mul2Context_delay_22_isFull <= SBox5Stage_mul2Context_delay_21_isFull;
    SBox5Stage_mul2Context_delay_22_fullRound <= SBox5Stage_mul2Context_delay_21_fullRound;
    SBox5Stage_mul2Context_delay_22_partialRound <= SBox5Stage_mul2Context_delay_21_partialRound;
    SBox5Stage_mul2Context_delay_22_stateIndex <= SBox5Stage_mul2Context_delay_21_stateIndex;
    SBox5Stage_mul2Context_delay_22_stateSize <= SBox5Stage_mul2Context_delay_21_stateSize;
    SBox5Stage_mul2Context_delay_22_stateID <= SBox5Stage_mul2Context_delay_21_stateID;
    SBox5Stage_mul2Context_delay_22_stateElements_0 <= SBox5Stage_mul2Context_delay_21_stateElements_0;
    SBox5Stage_mul2Context_delay_22_stateElements_1 <= SBox5Stage_mul2Context_delay_21_stateElements_1;
    SBox5Stage_mul2Context_delay_22_stateElements_2 <= SBox5Stage_mul2Context_delay_21_stateElements_2;
    SBox5Stage_mul2Context_delay_22_stateElements_3 <= SBox5Stage_mul2Context_delay_21_stateElements_3;
    SBox5Stage_mul2Context_delay_22_stateElements_4 <= SBox5Stage_mul2Context_delay_21_stateElements_4;
    SBox5Stage_mul2Context_delay_22_stateElements_5 <= SBox5Stage_mul2Context_delay_21_stateElements_5;
    SBox5Stage_mul2Context_delay_22_stateElements_6 <= SBox5Stage_mul2Context_delay_21_stateElements_6;
    SBox5Stage_mul2Context_delay_22_stateElements_7 <= SBox5Stage_mul2Context_delay_21_stateElements_7;
    SBox5Stage_mul2Context_delay_22_stateElements_8 <= SBox5Stage_mul2Context_delay_21_stateElements_8;
    SBox5Stage_mul2Context_delay_22_stateElements_9 <= SBox5Stage_mul2Context_delay_21_stateElements_9;
    SBox5Stage_mul2Context_delay_22_stateElements_10 <= SBox5Stage_mul2Context_delay_21_stateElements_10;
    SBox5Stage_mul2Context_delay_23_isFull <= SBox5Stage_mul2Context_delay_22_isFull;
    SBox5Stage_mul2Context_delay_23_fullRound <= SBox5Stage_mul2Context_delay_22_fullRound;
    SBox5Stage_mul2Context_delay_23_partialRound <= SBox5Stage_mul2Context_delay_22_partialRound;
    SBox5Stage_mul2Context_delay_23_stateIndex <= SBox5Stage_mul2Context_delay_22_stateIndex;
    SBox5Stage_mul2Context_delay_23_stateSize <= SBox5Stage_mul2Context_delay_22_stateSize;
    SBox5Stage_mul2Context_delay_23_stateID <= SBox5Stage_mul2Context_delay_22_stateID;
    SBox5Stage_mul2Context_delay_23_stateElements_0 <= SBox5Stage_mul2Context_delay_22_stateElements_0;
    SBox5Stage_mul2Context_delay_23_stateElements_1 <= SBox5Stage_mul2Context_delay_22_stateElements_1;
    SBox5Stage_mul2Context_delay_23_stateElements_2 <= SBox5Stage_mul2Context_delay_22_stateElements_2;
    SBox5Stage_mul2Context_delay_23_stateElements_3 <= SBox5Stage_mul2Context_delay_22_stateElements_3;
    SBox5Stage_mul2Context_delay_23_stateElements_4 <= SBox5Stage_mul2Context_delay_22_stateElements_4;
    SBox5Stage_mul2Context_delay_23_stateElements_5 <= SBox5Stage_mul2Context_delay_22_stateElements_5;
    SBox5Stage_mul2Context_delay_23_stateElements_6 <= SBox5Stage_mul2Context_delay_22_stateElements_6;
    SBox5Stage_mul2Context_delay_23_stateElements_7 <= SBox5Stage_mul2Context_delay_22_stateElements_7;
    SBox5Stage_mul2Context_delay_23_stateElements_8 <= SBox5Stage_mul2Context_delay_22_stateElements_8;
    SBox5Stage_mul2Context_delay_23_stateElements_9 <= SBox5Stage_mul2Context_delay_22_stateElements_9;
    SBox5Stage_mul2Context_delay_23_stateElements_10 <= SBox5Stage_mul2Context_delay_22_stateElements_10;
    SBox5Stage_mul2Context_delay_24_isFull <= SBox5Stage_mul2Context_delay_23_isFull;
    SBox5Stage_mul2Context_delay_24_fullRound <= SBox5Stage_mul2Context_delay_23_fullRound;
    SBox5Stage_mul2Context_delay_24_partialRound <= SBox5Stage_mul2Context_delay_23_partialRound;
    SBox5Stage_mul2Context_delay_24_stateIndex <= SBox5Stage_mul2Context_delay_23_stateIndex;
    SBox5Stage_mul2Context_delay_24_stateSize <= SBox5Stage_mul2Context_delay_23_stateSize;
    SBox5Stage_mul2Context_delay_24_stateID <= SBox5Stage_mul2Context_delay_23_stateID;
    SBox5Stage_mul2Context_delay_24_stateElements_0 <= SBox5Stage_mul2Context_delay_23_stateElements_0;
    SBox5Stage_mul2Context_delay_24_stateElements_1 <= SBox5Stage_mul2Context_delay_23_stateElements_1;
    SBox5Stage_mul2Context_delay_24_stateElements_2 <= SBox5Stage_mul2Context_delay_23_stateElements_2;
    SBox5Stage_mul2Context_delay_24_stateElements_3 <= SBox5Stage_mul2Context_delay_23_stateElements_3;
    SBox5Stage_mul2Context_delay_24_stateElements_4 <= SBox5Stage_mul2Context_delay_23_stateElements_4;
    SBox5Stage_mul2Context_delay_24_stateElements_5 <= SBox5Stage_mul2Context_delay_23_stateElements_5;
    SBox5Stage_mul2Context_delay_24_stateElements_6 <= SBox5Stage_mul2Context_delay_23_stateElements_6;
    SBox5Stage_mul2Context_delay_24_stateElements_7 <= SBox5Stage_mul2Context_delay_23_stateElements_7;
    SBox5Stage_mul2Context_delay_24_stateElements_8 <= SBox5Stage_mul2Context_delay_23_stateElements_8;
    SBox5Stage_mul2Context_delay_24_stateElements_9 <= SBox5Stage_mul2Context_delay_23_stateElements_9;
    SBox5Stage_mul2Context_delay_24_stateElements_10 <= SBox5Stage_mul2Context_delay_23_stateElements_10;
    SBox5Stage_mul2Context_delay_25_isFull <= SBox5Stage_mul2Context_delay_24_isFull;
    SBox5Stage_mul2Context_delay_25_fullRound <= SBox5Stage_mul2Context_delay_24_fullRound;
    SBox5Stage_mul2Context_delay_25_partialRound <= SBox5Stage_mul2Context_delay_24_partialRound;
    SBox5Stage_mul2Context_delay_25_stateIndex <= SBox5Stage_mul2Context_delay_24_stateIndex;
    SBox5Stage_mul2Context_delay_25_stateSize <= SBox5Stage_mul2Context_delay_24_stateSize;
    SBox5Stage_mul2Context_delay_25_stateID <= SBox5Stage_mul2Context_delay_24_stateID;
    SBox5Stage_mul2Context_delay_25_stateElements_0 <= SBox5Stage_mul2Context_delay_24_stateElements_0;
    SBox5Stage_mul2Context_delay_25_stateElements_1 <= SBox5Stage_mul2Context_delay_24_stateElements_1;
    SBox5Stage_mul2Context_delay_25_stateElements_2 <= SBox5Stage_mul2Context_delay_24_stateElements_2;
    SBox5Stage_mul2Context_delay_25_stateElements_3 <= SBox5Stage_mul2Context_delay_24_stateElements_3;
    SBox5Stage_mul2Context_delay_25_stateElements_4 <= SBox5Stage_mul2Context_delay_24_stateElements_4;
    SBox5Stage_mul2Context_delay_25_stateElements_5 <= SBox5Stage_mul2Context_delay_24_stateElements_5;
    SBox5Stage_mul2Context_delay_25_stateElements_6 <= SBox5Stage_mul2Context_delay_24_stateElements_6;
    SBox5Stage_mul2Context_delay_25_stateElements_7 <= SBox5Stage_mul2Context_delay_24_stateElements_7;
    SBox5Stage_mul2Context_delay_25_stateElements_8 <= SBox5Stage_mul2Context_delay_24_stateElements_8;
    SBox5Stage_mul2Context_delay_25_stateElements_9 <= SBox5Stage_mul2Context_delay_24_stateElements_9;
    SBox5Stage_mul2Context_delay_25_stateElements_10 <= SBox5Stage_mul2Context_delay_24_stateElements_10;
    SBox5Stage_mul2Context_delay_26_isFull <= SBox5Stage_mul2Context_delay_25_isFull;
    SBox5Stage_mul2Context_delay_26_fullRound <= SBox5Stage_mul2Context_delay_25_fullRound;
    SBox5Stage_mul2Context_delay_26_partialRound <= SBox5Stage_mul2Context_delay_25_partialRound;
    SBox5Stage_mul2Context_delay_26_stateIndex <= SBox5Stage_mul2Context_delay_25_stateIndex;
    SBox5Stage_mul2Context_delay_26_stateSize <= SBox5Stage_mul2Context_delay_25_stateSize;
    SBox5Stage_mul2Context_delay_26_stateID <= SBox5Stage_mul2Context_delay_25_stateID;
    SBox5Stage_mul2Context_delay_26_stateElements_0 <= SBox5Stage_mul2Context_delay_25_stateElements_0;
    SBox5Stage_mul2Context_delay_26_stateElements_1 <= SBox5Stage_mul2Context_delay_25_stateElements_1;
    SBox5Stage_mul2Context_delay_26_stateElements_2 <= SBox5Stage_mul2Context_delay_25_stateElements_2;
    SBox5Stage_mul2Context_delay_26_stateElements_3 <= SBox5Stage_mul2Context_delay_25_stateElements_3;
    SBox5Stage_mul2Context_delay_26_stateElements_4 <= SBox5Stage_mul2Context_delay_25_stateElements_4;
    SBox5Stage_mul2Context_delay_26_stateElements_5 <= SBox5Stage_mul2Context_delay_25_stateElements_5;
    SBox5Stage_mul2Context_delay_26_stateElements_6 <= SBox5Stage_mul2Context_delay_25_stateElements_6;
    SBox5Stage_mul2Context_delay_26_stateElements_7 <= SBox5Stage_mul2Context_delay_25_stateElements_7;
    SBox5Stage_mul2Context_delay_26_stateElements_8 <= SBox5Stage_mul2Context_delay_25_stateElements_8;
    SBox5Stage_mul2Context_delay_26_stateElements_9 <= SBox5Stage_mul2Context_delay_25_stateElements_9;
    SBox5Stage_mul2Context_delay_26_stateElements_10 <= SBox5Stage_mul2Context_delay_25_stateElements_10;
    SBox5Stage_mul2Context_delay_27_isFull <= SBox5Stage_mul2Context_delay_26_isFull;
    SBox5Stage_mul2Context_delay_27_fullRound <= SBox5Stage_mul2Context_delay_26_fullRound;
    SBox5Stage_mul2Context_delay_27_partialRound <= SBox5Stage_mul2Context_delay_26_partialRound;
    SBox5Stage_mul2Context_delay_27_stateIndex <= SBox5Stage_mul2Context_delay_26_stateIndex;
    SBox5Stage_mul2Context_delay_27_stateSize <= SBox5Stage_mul2Context_delay_26_stateSize;
    SBox5Stage_mul2Context_delay_27_stateID <= SBox5Stage_mul2Context_delay_26_stateID;
    SBox5Stage_mul2Context_delay_27_stateElements_0 <= SBox5Stage_mul2Context_delay_26_stateElements_0;
    SBox5Stage_mul2Context_delay_27_stateElements_1 <= SBox5Stage_mul2Context_delay_26_stateElements_1;
    SBox5Stage_mul2Context_delay_27_stateElements_2 <= SBox5Stage_mul2Context_delay_26_stateElements_2;
    SBox5Stage_mul2Context_delay_27_stateElements_3 <= SBox5Stage_mul2Context_delay_26_stateElements_3;
    SBox5Stage_mul2Context_delay_27_stateElements_4 <= SBox5Stage_mul2Context_delay_26_stateElements_4;
    SBox5Stage_mul2Context_delay_27_stateElements_5 <= SBox5Stage_mul2Context_delay_26_stateElements_5;
    SBox5Stage_mul2Context_delay_27_stateElements_6 <= SBox5Stage_mul2Context_delay_26_stateElements_6;
    SBox5Stage_mul2Context_delay_27_stateElements_7 <= SBox5Stage_mul2Context_delay_26_stateElements_7;
    SBox5Stage_mul2Context_delay_27_stateElements_8 <= SBox5Stage_mul2Context_delay_26_stateElements_8;
    SBox5Stage_mul2Context_delay_27_stateElements_9 <= SBox5Stage_mul2Context_delay_26_stateElements_9;
    SBox5Stage_mul2Context_delay_27_stateElements_10 <= SBox5Stage_mul2Context_delay_26_stateElements_10;
    SBox5Stage_mul2Context_delay_28_isFull <= SBox5Stage_mul2Context_delay_27_isFull;
    SBox5Stage_mul2Context_delay_28_fullRound <= SBox5Stage_mul2Context_delay_27_fullRound;
    SBox5Stage_mul2Context_delay_28_partialRound <= SBox5Stage_mul2Context_delay_27_partialRound;
    SBox5Stage_mul2Context_delay_28_stateIndex <= SBox5Stage_mul2Context_delay_27_stateIndex;
    SBox5Stage_mul2Context_delay_28_stateSize <= SBox5Stage_mul2Context_delay_27_stateSize;
    SBox5Stage_mul2Context_delay_28_stateID <= SBox5Stage_mul2Context_delay_27_stateID;
    SBox5Stage_mul2Context_delay_28_stateElements_0 <= SBox5Stage_mul2Context_delay_27_stateElements_0;
    SBox5Stage_mul2Context_delay_28_stateElements_1 <= SBox5Stage_mul2Context_delay_27_stateElements_1;
    SBox5Stage_mul2Context_delay_28_stateElements_2 <= SBox5Stage_mul2Context_delay_27_stateElements_2;
    SBox5Stage_mul2Context_delay_28_stateElements_3 <= SBox5Stage_mul2Context_delay_27_stateElements_3;
    SBox5Stage_mul2Context_delay_28_stateElements_4 <= SBox5Stage_mul2Context_delay_27_stateElements_4;
    SBox5Stage_mul2Context_delay_28_stateElements_5 <= SBox5Stage_mul2Context_delay_27_stateElements_5;
    SBox5Stage_mul2Context_delay_28_stateElements_6 <= SBox5Stage_mul2Context_delay_27_stateElements_6;
    SBox5Stage_mul2Context_delay_28_stateElements_7 <= SBox5Stage_mul2Context_delay_27_stateElements_7;
    SBox5Stage_mul2Context_delay_28_stateElements_8 <= SBox5Stage_mul2Context_delay_27_stateElements_8;
    SBox5Stage_mul2Context_delay_28_stateElements_9 <= SBox5Stage_mul2Context_delay_27_stateElements_9;
    SBox5Stage_mul2Context_delay_28_stateElements_10 <= SBox5Stage_mul2Context_delay_27_stateElements_10;
    SBox5Stage_mul2Context_delay_29_isFull <= SBox5Stage_mul2Context_delay_28_isFull;
    SBox5Stage_mul2Context_delay_29_fullRound <= SBox5Stage_mul2Context_delay_28_fullRound;
    SBox5Stage_mul2Context_delay_29_partialRound <= SBox5Stage_mul2Context_delay_28_partialRound;
    SBox5Stage_mul2Context_delay_29_stateIndex <= SBox5Stage_mul2Context_delay_28_stateIndex;
    SBox5Stage_mul2Context_delay_29_stateSize <= SBox5Stage_mul2Context_delay_28_stateSize;
    SBox5Stage_mul2Context_delay_29_stateID <= SBox5Stage_mul2Context_delay_28_stateID;
    SBox5Stage_mul2Context_delay_29_stateElements_0 <= SBox5Stage_mul2Context_delay_28_stateElements_0;
    SBox5Stage_mul2Context_delay_29_stateElements_1 <= SBox5Stage_mul2Context_delay_28_stateElements_1;
    SBox5Stage_mul2Context_delay_29_stateElements_2 <= SBox5Stage_mul2Context_delay_28_stateElements_2;
    SBox5Stage_mul2Context_delay_29_stateElements_3 <= SBox5Stage_mul2Context_delay_28_stateElements_3;
    SBox5Stage_mul2Context_delay_29_stateElements_4 <= SBox5Stage_mul2Context_delay_28_stateElements_4;
    SBox5Stage_mul2Context_delay_29_stateElements_5 <= SBox5Stage_mul2Context_delay_28_stateElements_5;
    SBox5Stage_mul2Context_delay_29_stateElements_6 <= SBox5Stage_mul2Context_delay_28_stateElements_6;
    SBox5Stage_mul2Context_delay_29_stateElements_7 <= SBox5Stage_mul2Context_delay_28_stateElements_7;
    SBox5Stage_mul2Context_delay_29_stateElements_8 <= SBox5Stage_mul2Context_delay_28_stateElements_8;
    SBox5Stage_mul2Context_delay_29_stateElements_9 <= SBox5Stage_mul2Context_delay_28_stateElements_9;
    SBox5Stage_mul2Context_delay_29_stateElements_10 <= SBox5Stage_mul2Context_delay_28_stateElements_10;
    SBox5Stage_mul2Context_delay_30_isFull <= SBox5Stage_mul2Context_delay_29_isFull;
    SBox5Stage_mul2Context_delay_30_fullRound <= SBox5Stage_mul2Context_delay_29_fullRound;
    SBox5Stage_mul2Context_delay_30_partialRound <= SBox5Stage_mul2Context_delay_29_partialRound;
    SBox5Stage_mul2Context_delay_30_stateIndex <= SBox5Stage_mul2Context_delay_29_stateIndex;
    SBox5Stage_mul2Context_delay_30_stateSize <= SBox5Stage_mul2Context_delay_29_stateSize;
    SBox5Stage_mul2Context_delay_30_stateID <= SBox5Stage_mul2Context_delay_29_stateID;
    SBox5Stage_mul2Context_delay_30_stateElements_0 <= SBox5Stage_mul2Context_delay_29_stateElements_0;
    SBox5Stage_mul2Context_delay_30_stateElements_1 <= SBox5Stage_mul2Context_delay_29_stateElements_1;
    SBox5Stage_mul2Context_delay_30_stateElements_2 <= SBox5Stage_mul2Context_delay_29_stateElements_2;
    SBox5Stage_mul2Context_delay_30_stateElements_3 <= SBox5Stage_mul2Context_delay_29_stateElements_3;
    SBox5Stage_mul2Context_delay_30_stateElements_4 <= SBox5Stage_mul2Context_delay_29_stateElements_4;
    SBox5Stage_mul2Context_delay_30_stateElements_5 <= SBox5Stage_mul2Context_delay_29_stateElements_5;
    SBox5Stage_mul2Context_delay_30_stateElements_6 <= SBox5Stage_mul2Context_delay_29_stateElements_6;
    SBox5Stage_mul2Context_delay_30_stateElements_7 <= SBox5Stage_mul2Context_delay_29_stateElements_7;
    SBox5Stage_mul2Context_delay_30_stateElements_8 <= SBox5Stage_mul2Context_delay_29_stateElements_8;
    SBox5Stage_mul2Context_delay_30_stateElements_9 <= SBox5Stage_mul2Context_delay_29_stateElements_9;
    SBox5Stage_mul2Context_delay_30_stateElements_10 <= SBox5Stage_mul2Context_delay_29_stateElements_10;
    SBox5Stage_mul2Context_delay_31_isFull <= SBox5Stage_mul2Context_delay_30_isFull;
    SBox5Stage_mul2Context_delay_31_fullRound <= SBox5Stage_mul2Context_delay_30_fullRound;
    SBox5Stage_mul2Context_delay_31_partialRound <= SBox5Stage_mul2Context_delay_30_partialRound;
    SBox5Stage_mul2Context_delay_31_stateIndex <= SBox5Stage_mul2Context_delay_30_stateIndex;
    SBox5Stage_mul2Context_delay_31_stateSize <= SBox5Stage_mul2Context_delay_30_stateSize;
    SBox5Stage_mul2Context_delay_31_stateID <= SBox5Stage_mul2Context_delay_30_stateID;
    SBox5Stage_mul2Context_delay_31_stateElements_0 <= SBox5Stage_mul2Context_delay_30_stateElements_0;
    SBox5Stage_mul2Context_delay_31_stateElements_1 <= SBox5Stage_mul2Context_delay_30_stateElements_1;
    SBox5Stage_mul2Context_delay_31_stateElements_2 <= SBox5Stage_mul2Context_delay_30_stateElements_2;
    SBox5Stage_mul2Context_delay_31_stateElements_3 <= SBox5Stage_mul2Context_delay_30_stateElements_3;
    SBox5Stage_mul2Context_delay_31_stateElements_4 <= SBox5Stage_mul2Context_delay_30_stateElements_4;
    SBox5Stage_mul2Context_delay_31_stateElements_5 <= SBox5Stage_mul2Context_delay_30_stateElements_5;
    SBox5Stage_mul2Context_delay_31_stateElements_6 <= SBox5Stage_mul2Context_delay_30_stateElements_6;
    SBox5Stage_mul2Context_delay_31_stateElements_7 <= SBox5Stage_mul2Context_delay_30_stateElements_7;
    SBox5Stage_mul2Context_delay_31_stateElements_8 <= SBox5Stage_mul2Context_delay_30_stateElements_8;
    SBox5Stage_mul2Context_delay_31_stateElements_9 <= SBox5Stage_mul2Context_delay_30_stateElements_9;
    SBox5Stage_mul2Context_delay_31_stateElements_10 <= SBox5Stage_mul2Context_delay_30_stateElements_10;
    SBox5Stage_mul2Context_delay_32_isFull <= SBox5Stage_mul2Context_delay_31_isFull;
    SBox5Stage_mul2Context_delay_32_fullRound <= SBox5Stage_mul2Context_delay_31_fullRound;
    SBox5Stage_mul2Context_delay_32_partialRound <= SBox5Stage_mul2Context_delay_31_partialRound;
    SBox5Stage_mul2Context_delay_32_stateIndex <= SBox5Stage_mul2Context_delay_31_stateIndex;
    SBox5Stage_mul2Context_delay_32_stateSize <= SBox5Stage_mul2Context_delay_31_stateSize;
    SBox5Stage_mul2Context_delay_32_stateID <= SBox5Stage_mul2Context_delay_31_stateID;
    SBox5Stage_mul2Context_delay_32_stateElements_0 <= SBox5Stage_mul2Context_delay_31_stateElements_0;
    SBox5Stage_mul2Context_delay_32_stateElements_1 <= SBox5Stage_mul2Context_delay_31_stateElements_1;
    SBox5Stage_mul2Context_delay_32_stateElements_2 <= SBox5Stage_mul2Context_delay_31_stateElements_2;
    SBox5Stage_mul2Context_delay_32_stateElements_3 <= SBox5Stage_mul2Context_delay_31_stateElements_3;
    SBox5Stage_mul2Context_delay_32_stateElements_4 <= SBox5Stage_mul2Context_delay_31_stateElements_4;
    SBox5Stage_mul2Context_delay_32_stateElements_5 <= SBox5Stage_mul2Context_delay_31_stateElements_5;
    SBox5Stage_mul2Context_delay_32_stateElements_6 <= SBox5Stage_mul2Context_delay_31_stateElements_6;
    SBox5Stage_mul2Context_delay_32_stateElements_7 <= SBox5Stage_mul2Context_delay_31_stateElements_7;
    SBox5Stage_mul2Context_delay_32_stateElements_8 <= SBox5Stage_mul2Context_delay_31_stateElements_8;
    SBox5Stage_mul2Context_delay_32_stateElements_9 <= SBox5Stage_mul2Context_delay_31_stateElements_9;
    SBox5Stage_mul2Context_delay_32_stateElements_10 <= SBox5Stage_mul2Context_delay_31_stateElements_10;
    SBox5Stage_mul2Context_delay_33_isFull <= SBox5Stage_mul2Context_delay_32_isFull;
    SBox5Stage_mul2Context_delay_33_fullRound <= SBox5Stage_mul2Context_delay_32_fullRound;
    SBox5Stage_mul2Context_delay_33_partialRound <= SBox5Stage_mul2Context_delay_32_partialRound;
    SBox5Stage_mul2Context_delay_33_stateIndex <= SBox5Stage_mul2Context_delay_32_stateIndex;
    SBox5Stage_mul2Context_delay_33_stateSize <= SBox5Stage_mul2Context_delay_32_stateSize;
    SBox5Stage_mul2Context_delay_33_stateID <= SBox5Stage_mul2Context_delay_32_stateID;
    SBox5Stage_mul2Context_delay_33_stateElements_0 <= SBox5Stage_mul2Context_delay_32_stateElements_0;
    SBox5Stage_mul2Context_delay_33_stateElements_1 <= SBox5Stage_mul2Context_delay_32_stateElements_1;
    SBox5Stage_mul2Context_delay_33_stateElements_2 <= SBox5Stage_mul2Context_delay_32_stateElements_2;
    SBox5Stage_mul2Context_delay_33_stateElements_3 <= SBox5Stage_mul2Context_delay_32_stateElements_3;
    SBox5Stage_mul2Context_delay_33_stateElements_4 <= SBox5Stage_mul2Context_delay_32_stateElements_4;
    SBox5Stage_mul2Context_delay_33_stateElements_5 <= SBox5Stage_mul2Context_delay_32_stateElements_5;
    SBox5Stage_mul2Context_delay_33_stateElements_6 <= SBox5Stage_mul2Context_delay_32_stateElements_6;
    SBox5Stage_mul2Context_delay_33_stateElements_7 <= SBox5Stage_mul2Context_delay_32_stateElements_7;
    SBox5Stage_mul2Context_delay_33_stateElements_8 <= SBox5Stage_mul2Context_delay_32_stateElements_8;
    SBox5Stage_mul2Context_delay_33_stateElements_9 <= SBox5Stage_mul2Context_delay_32_stateElements_9;
    SBox5Stage_mul2Context_delay_33_stateElements_10 <= SBox5Stage_mul2Context_delay_32_stateElements_10;
    SBox5Stage_mul2Context_delay_34_isFull <= SBox5Stage_mul2Context_delay_33_isFull;
    SBox5Stage_mul2Context_delay_34_fullRound <= SBox5Stage_mul2Context_delay_33_fullRound;
    SBox5Stage_mul2Context_delay_34_partialRound <= SBox5Stage_mul2Context_delay_33_partialRound;
    SBox5Stage_mul2Context_delay_34_stateIndex <= SBox5Stage_mul2Context_delay_33_stateIndex;
    SBox5Stage_mul2Context_delay_34_stateSize <= SBox5Stage_mul2Context_delay_33_stateSize;
    SBox5Stage_mul2Context_delay_34_stateID <= SBox5Stage_mul2Context_delay_33_stateID;
    SBox5Stage_mul2Context_delay_34_stateElements_0 <= SBox5Stage_mul2Context_delay_33_stateElements_0;
    SBox5Stage_mul2Context_delay_34_stateElements_1 <= SBox5Stage_mul2Context_delay_33_stateElements_1;
    SBox5Stage_mul2Context_delay_34_stateElements_2 <= SBox5Stage_mul2Context_delay_33_stateElements_2;
    SBox5Stage_mul2Context_delay_34_stateElements_3 <= SBox5Stage_mul2Context_delay_33_stateElements_3;
    SBox5Stage_mul2Context_delay_34_stateElements_4 <= SBox5Stage_mul2Context_delay_33_stateElements_4;
    SBox5Stage_mul2Context_delay_34_stateElements_5 <= SBox5Stage_mul2Context_delay_33_stateElements_5;
    SBox5Stage_mul2Context_delay_34_stateElements_6 <= SBox5Stage_mul2Context_delay_33_stateElements_6;
    SBox5Stage_mul2Context_delay_34_stateElements_7 <= SBox5Stage_mul2Context_delay_33_stateElements_7;
    SBox5Stage_mul2Context_delay_34_stateElements_8 <= SBox5Stage_mul2Context_delay_33_stateElements_8;
    SBox5Stage_mul2Context_delay_34_stateElements_9 <= SBox5Stage_mul2Context_delay_33_stateElements_9;
    SBox5Stage_mul2Context_delay_34_stateElements_10 <= SBox5Stage_mul2Context_delay_33_stateElements_10;
    SBox5Stage_mul2Context_delay_35_isFull <= SBox5Stage_mul2Context_delay_34_isFull;
    SBox5Stage_mul2Context_delay_35_fullRound <= SBox5Stage_mul2Context_delay_34_fullRound;
    SBox5Stage_mul2Context_delay_35_partialRound <= SBox5Stage_mul2Context_delay_34_partialRound;
    SBox5Stage_mul2Context_delay_35_stateIndex <= SBox5Stage_mul2Context_delay_34_stateIndex;
    SBox5Stage_mul2Context_delay_35_stateSize <= SBox5Stage_mul2Context_delay_34_stateSize;
    SBox5Stage_mul2Context_delay_35_stateID <= SBox5Stage_mul2Context_delay_34_stateID;
    SBox5Stage_mul2Context_delay_35_stateElements_0 <= SBox5Stage_mul2Context_delay_34_stateElements_0;
    SBox5Stage_mul2Context_delay_35_stateElements_1 <= SBox5Stage_mul2Context_delay_34_stateElements_1;
    SBox5Stage_mul2Context_delay_35_stateElements_2 <= SBox5Stage_mul2Context_delay_34_stateElements_2;
    SBox5Stage_mul2Context_delay_35_stateElements_3 <= SBox5Stage_mul2Context_delay_34_stateElements_3;
    SBox5Stage_mul2Context_delay_35_stateElements_4 <= SBox5Stage_mul2Context_delay_34_stateElements_4;
    SBox5Stage_mul2Context_delay_35_stateElements_5 <= SBox5Stage_mul2Context_delay_34_stateElements_5;
    SBox5Stage_mul2Context_delay_35_stateElements_6 <= SBox5Stage_mul2Context_delay_34_stateElements_6;
    SBox5Stage_mul2Context_delay_35_stateElements_7 <= SBox5Stage_mul2Context_delay_34_stateElements_7;
    SBox5Stage_mul2Context_delay_35_stateElements_8 <= SBox5Stage_mul2Context_delay_34_stateElements_8;
    SBox5Stage_mul2Context_delay_35_stateElements_9 <= SBox5Stage_mul2Context_delay_34_stateElements_9;
    SBox5Stage_mul2Context_delay_35_stateElements_10 <= SBox5Stage_mul2Context_delay_34_stateElements_10;
    SBox5Stage_mul2Context_delay_36_isFull <= SBox5Stage_mul2Context_delay_35_isFull;
    SBox5Stage_mul2Context_delay_36_fullRound <= SBox5Stage_mul2Context_delay_35_fullRound;
    SBox5Stage_mul2Context_delay_36_partialRound <= SBox5Stage_mul2Context_delay_35_partialRound;
    SBox5Stage_mul2Context_delay_36_stateIndex <= SBox5Stage_mul2Context_delay_35_stateIndex;
    SBox5Stage_mul2Context_delay_36_stateSize <= SBox5Stage_mul2Context_delay_35_stateSize;
    SBox5Stage_mul2Context_delay_36_stateID <= SBox5Stage_mul2Context_delay_35_stateID;
    SBox5Stage_mul2Context_delay_36_stateElements_0 <= SBox5Stage_mul2Context_delay_35_stateElements_0;
    SBox5Stage_mul2Context_delay_36_stateElements_1 <= SBox5Stage_mul2Context_delay_35_stateElements_1;
    SBox5Stage_mul2Context_delay_36_stateElements_2 <= SBox5Stage_mul2Context_delay_35_stateElements_2;
    SBox5Stage_mul2Context_delay_36_stateElements_3 <= SBox5Stage_mul2Context_delay_35_stateElements_3;
    SBox5Stage_mul2Context_delay_36_stateElements_4 <= SBox5Stage_mul2Context_delay_35_stateElements_4;
    SBox5Stage_mul2Context_delay_36_stateElements_5 <= SBox5Stage_mul2Context_delay_35_stateElements_5;
    SBox5Stage_mul2Context_delay_36_stateElements_6 <= SBox5Stage_mul2Context_delay_35_stateElements_6;
    SBox5Stage_mul2Context_delay_36_stateElements_7 <= SBox5Stage_mul2Context_delay_35_stateElements_7;
    SBox5Stage_mul2Context_delay_36_stateElements_8 <= SBox5Stage_mul2Context_delay_35_stateElements_8;
    SBox5Stage_mul2Context_delay_36_stateElements_9 <= SBox5Stage_mul2Context_delay_35_stateElements_9;
    SBox5Stage_mul2Context_delay_36_stateElements_10 <= SBox5Stage_mul2Context_delay_35_stateElements_10;
    SBox5Stage_mul2Context_delay_37_isFull <= SBox5Stage_mul2Context_delay_36_isFull;
    SBox5Stage_mul2Context_delay_37_fullRound <= SBox5Stage_mul2Context_delay_36_fullRound;
    SBox5Stage_mul2Context_delay_37_partialRound <= SBox5Stage_mul2Context_delay_36_partialRound;
    SBox5Stage_mul2Context_delay_37_stateIndex <= SBox5Stage_mul2Context_delay_36_stateIndex;
    SBox5Stage_mul2Context_delay_37_stateSize <= SBox5Stage_mul2Context_delay_36_stateSize;
    SBox5Stage_mul2Context_delay_37_stateID <= SBox5Stage_mul2Context_delay_36_stateID;
    SBox5Stage_mul2Context_delay_37_stateElements_0 <= SBox5Stage_mul2Context_delay_36_stateElements_0;
    SBox5Stage_mul2Context_delay_37_stateElements_1 <= SBox5Stage_mul2Context_delay_36_stateElements_1;
    SBox5Stage_mul2Context_delay_37_stateElements_2 <= SBox5Stage_mul2Context_delay_36_stateElements_2;
    SBox5Stage_mul2Context_delay_37_stateElements_3 <= SBox5Stage_mul2Context_delay_36_stateElements_3;
    SBox5Stage_mul2Context_delay_37_stateElements_4 <= SBox5Stage_mul2Context_delay_36_stateElements_4;
    SBox5Stage_mul2Context_delay_37_stateElements_5 <= SBox5Stage_mul2Context_delay_36_stateElements_5;
    SBox5Stage_mul2Context_delay_37_stateElements_6 <= SBox5Stage_mul2Context_delay_36_stateElements_6;
    SBox5Stage_mul2Context_delay_37_stateElements_7 <= SBox5Stage_mul2Context_delay_36_stateElements_7;
    SBox5Stage_mul2Context_delay_37_stateElements_8 <= SBox5Stage_mul2Context_delay_36_stateElements_8;
    SBox5Stage_mul2Context_delay_37_stateElements_9 <= SBox5Stage_mul2Context_delay_36_stateElements_9;
    SBox5Stage_mul2Context_delay_37_stateElements_10 <= SBox5Stage_mul2Context_delay_36_stateElements_10;
    SBox5Stage_mul2Context_delay_38_isFull <= SBox5Stage_mul2Context_delay_37_isFull;
    SBox5Stage_mul2Context_delay_38_fullRound <= SBox5Stage_mul2Context_delay_37_fullRound;
    SBox5Stage_mul2Context_delay_38_partialRound <= SBox5Stage_mul2Context_delay_37_partialRound;
    SBox5Stage_mul2Context_delay_38_stateIndex <= SBox5Stage_mul2Context_delay_37_stateIndex;
    SBox5Stage_mul2Context_delay_38_stateSize <= SBox5Stage_mul2Context_delay_37_stateSize;
    SBox5Stage_mul2Context_delay_38_stateID <= SBox5Stage_mul2Context_delay_37_stateID;
    SBox5Stage_mul2Context_delay_38_stateElements_0 <= SBox5Stage_mul2Context_delay_37_stateElements_0;
    SBox5Stage_mul2Context_delay_38_stateElements_1 <= SBox5Stage_mul2Context_delay_37_stateElements_1;
    SBox5Stage_mul2Context_delay_38_stateElements_2 <= SBox5Stage_mul2Context_delay_37_stateElements_2;
    SBox5Stage_mul2Context_delay_38_stateElements_3 <= SBox5Stage_mul2Context_delay_37_stateElements_3;
    SBox5Stage_mul2Context_delay_38_stateElements_4 <= SBox5Stage_mul2Context_delay_37_stateElements_4;
    SBox5Stage_mul2Context_delay_38_stateElements_5 <= SBox5Stage_mul2Context_delay_37_stateElements_5;
    SBox5Stage_mul2Context_delay_38_stateElements_6 <= SBox5Stage_mul2Context_delay_37_stateElements_6;
    SBox5Stage_mul2Context_delay_38_stateElements_7 <= SBox5Stage_mul2Context_delay_37_stateElements_7;
    SBox5Stage_mul2Context_delay_38_stateElements_8 <= SBox5Stage_mul2Context_delay_37_stateElements_8;
    SBox5Stage_mul2Context_delay_38_stateElements_9 <= SBox5Stage_mul2Context_delay_37_stateElements_9;
    SBox5Stage_mul2Context_delay_38_stateElements_10 <= SBox5Stage_mul2Context_delay_37_stateElements_10;
    SBox5Stage_mul2Context_delay_39_isFull <= SBox5Stage_mul2Context_delay_38_isFull;
    SBox5Stage_mul2Context_delay_39_fullRound <= SBox5Stage_mul2Context_delay_38_fullRound;
    SBox5Stage_mul2Context_delay_39_partialRound <= SBox5Stage_mul2Context_delay_38_partialRound;
    SBox5Stage_mul2Context_delay_39_stateIndex <= SBox5Stage_mul2Context_delay_38_stateIndex;
    SBox5Stage_mul2Context_delay_39_stateSize <= SBox5Stage_mul2Context_delay_38_stateSize;
    SBox5Stage_mul2Context_delay_39_stateID <= SBox5Stage_mul2Context_delay_38_stateID;
    SBox5Stage_mul2Context_delay_39_stateElements_0 <= SBox5Stage_mul2Context_delay_38_stateElements_0;
    SBox5Stage_mul2Context_delay_39_stateElements_1 <= SBox5Stage_mul2Context_delay_38_stateElements_1;
    SBox5Stage_mul2Context_delay_39_stateElements_2 <= SBox5Stage_mul2Context_delay_38_stateElements_2;
    SBox5Stage_mul2Context_delay_39_stateElements_3 <= SBox5Stage_mul2Context_delay_38_stateElements_3;
    SBox5Stage_mul2Context_delay_39_stateElements_4 <= SBox5Stage_mul2Context_delay_38_stateElements_4;
    SBox5Stage_mul2Context_delay_39_stateElements_5 <= SBox5Stage_mul2Context_delay_38_stateElements_5;
    SBox5Stage_mul2Context_delay_39_stateElements_6 <= SBox5Stage_mul2Context_delay_38_stateElements_6;
    SBox5Stage_mul2Context_delay_39_stateElements_7 <= SBox5Stage_mul2Context_delay_38_stateElements_7;
    SBox5Stage_mul2Context_delay_39_stateElements_8 <= SBox5Stage_mul2Context_delay_38_stateElements_8;
    SBox5Stage_mul2Context_delay_39_stateElements_9 <= SBox5Stage_mul2Context_delay_38_stateElements_9;
    SBox5Stage_mul2Context_delay_39_stateElements_10 <= SBox5Stage_mul2Context_delay_38_stateElements_10;
    SBox5Stage_mul2Context_delay_40_isFull <= SBox5Stage_mul2Context_delay_39_isFull;
    SBox5Stage_mul2Context_delay_40_fullRound <= SBox5Stage_mul2Context_delay_39_fullRound;
    SBox5Stage_mul2Context_delay_40_partialRound <= SBox5Stage_mul2Context_delay_39_partialRound;
    SBox5Stage_mul2Context_delay_40_stateIndex <= SBox5Stage_mul2Context_delay_39_stateIndex;
    SBox5Stage_mul2Context_delay_40_stateSize <= SBox5Stage_mul2Context_delay_39_stateSize;
    SBox5Stage_mul2Context_delay_40_stateID <= SBox5Stage_mul2Context_delay_39_stateID;
    SBox5Stage_mul2Context_delay_40_stateElements_0 <= SBox5Stage_mul2Context_delay_39_stateElements_0;
    SBox5Stage_mul2Context_delay_40_stateElements_1 <= SBox5Stage_mul2Context_delay_39_stateElements_1;
    SBox5Stage_mul2Context_delay_40_stateElements_2 <= SBox5Stage_mul2Context_delay_39_stateElements_2;
    SBox5Stage_mul2Context_delay_40_stateElements_3 <= SBox5Stage_mul2Context_delay_39_stateElements_3;
    SBox5Stage_mul2Context_delay_40_stateElements_4 <= SBox5Stage_mul2Context_delay_39_stateElements_4;
    SBox5Stage_mul2Context_delay_40_stateElements_5 <= SBox5Stage_mul2Context_delay_39_stateElements_5;
    SBox5Stage_mul2Context_delay_40_stateElements_6 <= SBox5Stage_mul2Context_delay_39_stateElements_6;
    SBox5Stage_mul2Context_delay_40_stateElements_7 <= SBox5Stage_mul2Context_delay_39_stateElements_7;
    SBox5Stage_mul2Context_delay_40_stateElements_8 <= SBox5Stage_mul2Context_delay_39_stateElements_8;
    SBox5Stage_mul2Context_delay_40_stateElements_9 <= SBox5Stage_mul2Context_delay_39_stateElements_9;
    SBox5Stage_mul2Context_delay_40_stateElements_10 <= SBox5Stage_mul2Context_delay_39_stateElements_10;
    SBox5Stage_mul2Context_delay_41_isFull <= SBox5Stage_mul2Context_delay_40_isFull;
    SBox5Stage_mul2Context_delay_41_fullRound <= SBox5Stage_mul2Context_delay_40_fullRound;
    SBox5Stage_mul2Context_delay_41_partialRound <= SBox5Stage_mul2Context_delay_40_partialRound;
    SBox5Stage_mul2Context_delay_41_stateIndex <= SBox5Stage_mul2Context_delay_40_stateIndex;
    SBox5Stage_mul2Context_delay_41_stateSize <= SBox5Stage_mul2Context_delay_40_stateSize;
    SBox5Stage_mul2Context_delay_41_stateID <= SBox5Stage_mul2Context_delay_40_stateID;
    SBox5Stage_mul2Context_delay_41_stateElements_0 <= SBox5Stage_mul2Context_delay_40_stateElements_0;
    SBox5Stage_mul2Context_delay_41_stateElements_1 <= SBox5Stage_mul2Context_delay_40_stateElements_1;
    SBox5Stage_mul2Context_delay_41_stateElements_2 <= SBox5Stage_mul2Context_delay_40_stateElements_2;
    SBox5Stage_mul2Context_delay_41_stateElements_3 <= SBox5Stage_mul2Context_delay_40_stateElements_3;
    SBox5Stage_mul2Context_delay_41_stateElements_4 <= SBox5Stage_mul2Context_delay_40_stateElements_4;
    SBox5Stage_mul2Context_delay_41_stateElements_5 <= SBox5Stage_mul2Context_delay_40_stateElements_5;
    SBox5Stage_mul2Context_delay_41_stateElements_6 <= SBox5Stage_mul2Context_delay_40_stateElements_6;
    SBox5Stage_mul2Context_delay_41_stateElements_7 <= SBox5Stage_mul2Context_delay_40_stateElements_7;
    SBox5Stage_mul2Context_delay_41_stateElements_8 <= SBox5Stage_mul2Context_delay_40_stateElements_8;
    SBox5Stage_mul2Context_delay_41_stateElements_9 <= SBox5Stage_mul2Context_delay_40_stateElements_9;
    SBox5Stage_mul2Context_delay_41_stateElements_10 <= SBox5Stage_mul2Context_delay_40_stateElements_10;
    SBox5Stage_mul2Context_delay_42_isFull <= SBox5Stage_mul2Context_delay_41_isFull;
    SBox5Stage_mul2Context_delay_42_fullRound <= SBox5Stage_mul2Context_delay_41_fullRound;
    SBox5Stage_mul2Context_delay_42_partialRound <= SBox5Stage_mul2Context_delay_41_partialRound;
    SBox5Stage_mul2Context_delay_42_stateIndex <= SBox5Stage_mul2Context_delay_41_stateIndex;
    SBox5Stage_mul2Context_delay_42_stateSize <= SBox5Stage_mul2Context_delay_41_stateSize;
    SBox5Stage_mul2Context_delay_42_stateID <= SBox5Stage_mul2Context_delay_41_stateID;
    SBox5Stage_mul2Context_delay_42_stateElements_0 <= SBox5Stage_mul2Context_delay_41_stateElements_0;
    SBox5Stage_mul2Context_delay_42_stateElements_1 <= SBox5Stage_mul2Context_delay_41_stateElements_1;
    SBox5Stage_mul2Context_delay_42_stateElements_2 <= SBox5Stage_mul2Context_delay_41_stateElements_2;
    SBox5Stage_mul2Context_delay_42_stateElements_3 <= SBox5Stage_mul2Context_delay_41_stateElements_3;
    SBox5Stage_mul2Context_delay_42_stateElements_4 <= SBox5Stage_mul2Context_delay_41_stateElements_4;
    SBox5Stage_mul2Context_delay_42_stateElements_5 <= SBox5Stage_mul2Context_delay_41_stateElements_5;
    SBox5Stage_mul2Context_delay_42_stateElements_6 <= SBox5Stage_mul2Context_delay_41_stateElements_6;
    SBox5Stage_mul2Context_delay_42_stateElements_7 <= SBox5Stage_mul2Context_delay_41_stateElements_7;
    SBox5Stage_mul2Context_delay_42_stateElements_8 <= SBox5Stage_mul2Context_delay_41_stateElements_8;
    SBox5Stage_mul2Context_delay_42_stateElements_9 <= SBox5Stage_mul2Context_delay_41_stateElements_9;
    SBox5Stage_mul2Context_delay_42_stateElements_10 <= SBox5Stage_mul2Context_delay_41_stateElements_10;
    SBox5Stage_mul2Context_delay_43_isFull <= SBox5Stage_mul2Context_delay_42_isFull;
    SBox5Stage_mul2Context_delay_43_fullRound <= SBox5Stage_mul2Context_delay_42_fullRound;
    SBox5Stage_mul2Context_delay_43_partialRound <= SBox5Stage_mul2Context_delay_42_partialRound;
    SBox5Stage_mul2Context_delay_43_stateIndex <= SBox5Stage_mul2Context_delay_42_stateIndex;
    SBox5Stage_mul2Context_delay_43_stateSize <= SBox5Stage_mul2Context_delay_42_stateSize;
    SBox5Stage_mul2Context_delay_43_stateID <= SBox5Stage_mul2Context_delay_42_stateID;
    SBox5Stage_mul2Context_delay_43_stateElements_0 <= SBox5Stage_mul2Context_delay_42_stateElements_0;
    SBox5Stage_mul2Context_delay_43_stateElements_1 <= SBox5Stage_mul2Context_delay_42_stateElements_1;
    SBox5Stage_mul2Context_delay_43_stateElements_2 <= SBox5Stage_mul2Context_delay_42_stateElements_2;
    SBox5Stage_mul2Context_delay_43_stateElements_3 <= SBox5Stage_mul2Context_delay_42_stateElements_3;
    SBox5Stage_mul2Context_delay_43_stateElements_4 <= SBox5Stage_mul2Context_delay_42_stateElements_4;
    SBox5Stage_mul2Context_delay_43_stateElements_5 <= SBox5Stage_mul2Context_delay_42_stateElements_5;
    SBox5Stage_mul2Context_delay_43_stateElements_6 <= SBox5Stage_mul2Context_delay_42_stateElements_6;
    SBox5Stage_mul2Context_delay_43_stateElements_7 <= SBox5Stage_mul2Context_delay_42_stateElements_7;
    SBox5Stage_mul2Context_delay_43_stateElements_8 <= SBox5Stage_mul2Context_delay_42_stateElements_8;
    SBox5Stage_mul2Context_delay_43_stateElements_9 <= SBox5Stage_mul2Context_delay_42_stateElements_9;
    SBox5Stage_mul2Context_delay_43_stateElements_10 <= SBox5Stage_mul2Context_delay_42_stateElements_10;
    SBox5Stage_mul2Context_delay_44_isFull <= SBox5Stage_mul2Context_delay_43_isFull;
    SBox5Stage_mul2Context_delay_44_fullRound <= SBox5Stage_mul2Context_delay_43_fullRound;
    SBox5Stage_mul2Context_delay_44_partialRound <= SBox5Stage_mul2Context_delay_43_partialRound;
    SBox5Stage_mul2Context_delay_44_stateIndex <= SBox5Stage_mul2Context_delay_43_stateIndex;
    SBox5Stage_mul2Context_delay_44_stateSize <= SBox5Stage_mul2Context_delay_43_stateSize;
    SBox5Stage_mul2Context_delay_44_stateID <= SBox5Stage_mul2Context_delay_43_stateID;
    SBox5Stage_mul2Context_delay_44_stateElements_0 <= SBox5Stage_mul2Context_delay_43_stateElements_0;
    SBox5Stage_mul2Context_delay_44_stateElements_1 <= SBox5Stage_mul2Context_delay_43_stateElements_1;
    SBox5Stage_mul2Context_delay_44_stateElements_2 <= SBox5Stage_mul2Context_delay_43_stateElements_2;
    SBox5Stage_mul2Context_delay_44_stateElements_3 <= SBox5Stage_mul2Context_delay_43_stateElements_3;
    SBox5Stage_mul2Context_delay_44_stateElements_4 <= SBox5Stage_mul2Context_delay_43_stateElements_4;
    SBox5Stage_mul2Context_delay_44_stateElements_5 <= SBox5Stage_mul2Context_delay_43_stateElements_5;
    SBox5Stage_mul2Context_delay_44_stateElements_6 <= SBox5Stage_mul2Context_delay_43_stateElements_6;
    SBox5Stage_mul2Context_delay_44_stateElements_7 <= SBox5Stage_mul2Context_delay_43_stateElements_7;
    SBox5Stage_mul2Context_delay_44_stateElements_8 <= SBox5Stage_mul2Context_delay_43_stateElements_8;
    SBox5Stage_mul2Context_delay_44_stateElements_9 <= SBox5Stage_mul2Context_delay_43_stateElements_9;
    SBox5Stage_mul2Context_delay_44_stateElements_10 <= SBox5Stage_mul2Context_delay_43_stateElements_10;
    SBox5Stage_mul2Context_delay_45_isFull <= SBox5Stage_mul2Context_delay_44_isFull;
    SBox5Stage_mul2Context_delay_45_fullRound <= SBox5Stage_mul2Context_delay_44_fullRound;
    SBox5Stage_mul2Context_delay_45_partialRound <= SBox5Stage_mul2Context_delay_44_partialRound;
    SBox5Stage_mul2Context_delay_45_stateIndex <= SBox5Stage_mul2Context_delay_44_stateIndex;
    SBox5Stage_mul2Context_delay_45_stateSize <= SBox5Stage_mul2Context_delay_44_stateSize;
    SBox5Stage_mul2Context_delay_45_stateID <= SBox5Stage_mul2Context_delay_44_stateID;
    SBox5Stage_mul2Context_delay_45_stateElements_0 <= SBox5Stage_mul2Context_delay_44_stateElements_0;
    SBox5Stage_mul2Context_delay_45_stateElements_1 <= SBox5Stage_mul2Context_delay_44_stateElements_1;
    SBox5Stage_mul2Context_delay_45_stateElements_2 <= SBox5Stage_mul2Context_delay_44_stateElements_2;
    SBox5Stage_mul2Context_delay_45_stateElements_3 <= SBox5Stage_mul2Context_delay_44_stateElements_3;
    SBox5Stage_mul2Context_delay_45_stateElements_4 <= SBox5Stage_mul2Context_delay_44_stateElements_4;
    SBox5Stage_mul2Context_delay_45_stateElements_5 <= SBox5Stage_mul2Context_delay_44_stateElements_5;
    SBox5Stage_mul2Context_delay_45_stateElements_6 <= SBox5Stage_mul2Context_delay_44_stateElements_6;
    SBox5Stage_mul2Context_delay_45_stateElements_7 <= SBox5Stage_mul2Context_delay_44_stateElements_7;
    SBox5Stage_mul2Context_delay_45_stateElements_8 <= SBox5Stage_mul2Context_delay_44_stateElements_8;
    SBox5Stage_mul2Context_delay_45_stateElements_9 <= SBox5Stage_mul2Context_delay_44_stateElements_9;
    SBox5Stage_mul2Context_delay_45_stateElements_10 <= SBox5Stage_mul2Context_delay_44_stateElements_10;
    SBox5Stage_mul2Context_delay_46_isFull <= SBox5Stage_mul2Context_delay_45_isFull;
    SBox5Stage_mul2Context_delay_46_fullRound <= SBox5Stage_mul2Context_delay_45_fullRound;
    SBox5Stage_mul2Context_delay_46_partialRound <= SBox5Stage_mul2Context_delay_45_partialRound;
    SBox5Stage_mul2Context_delay_46_stateIndex <= SBox5Stage_mul2Context_delay_45_stateIndex;
    SBox5Stage_mul2Context_delay_46_stateSize <= SBox5Stage_mul2Context_delay_45_stateSize;
    SBox5Stage_mul2Context_delay_46_stateID <= SBox5Stage_mul2Context_delay_45_stateID;
    SBox5Stage_mul2Context_delay_46_stateElements_0 <= SBox5Stage_mul2Context_delay_45_stateElements_0;
    SBox5Stage_mul2Context_delay_46_stateElements_1 <= SBox5Stage_mul2Context_delay_45_stateElements_1;
    SBox5Stage_mul2Context_delay_46_stateElements_2 <= SBox5Stage_mul2Context_delay_45_stateElements_2;
    SBox5Stage_mul2Context_delay_46_stateElements_3 <= SBox5Stage_mul2Context_delay_45_stateElements_3;
    SBox5Stage_mul2Context_delay_46_stateElements_4 <= SBox5Stage_mul2Context_delay_45_stateElements_4;
    SBox5Stage_mul2Context_delay_46_stateElements_5 <= SBox5Stage_mul2Context_delay_45_stateElements_5;
    SBox5Stage_mul2Context_delay_46_stateElements_6 <= SBox5Stage_mul2Context_delay_45_stateElements_6;
    SBox5Stage_mul2Context_delay_46_stateElements_7 <= SBox5Stage_mul2Context_delay_45_stateElements_7;
    SBox5Stage_mul2Context_delay_46_stateElements_8 <= SBox5Stage_mul2Context_delay_45_stateElements_8;
    SBox5Stage_mul2Context_delay_46_stateElements_9 <= SBox5Stage_mul2Context_delay_45_stateElements_9;
    SBox5Stage_mul2Context_delay_46_stateElements_10 <= SBox5Stage_mul2Context_delay_45_stateElements_10;
    SBox5Stage_mul2Context_delay_47_isFull <= SBox5Stage_mul2Context_delay_46_isFull;
    SBox5Stage_mul2Context_delay_47_fullRound <= SBox5Stage_mul2Context_delay_46_fullRound;
    SBox5Stage_mul2Context_delay_47_partialRound <= SBox5Stage_mul2Context_delay_46_partialRound;
    SBox5Stage_mul2Context_delay_47_stateIndex <= SBox5Stage_mul2Context_delay_46_stateIndex;
    SBox5Stage_mul2Context_delay_47_stateSize <= SBox5Stage_mul2Context_delay_46_stateSize;
    SBox5Stage_mul2Context_delay_47_stateID <= SBox5Stage_mul2Context_delay_46_stateID;
    SBox5Stage_mul2Context_delay_47_stateElements_0 <= SBox5Stage_mul2Context_delay_46_stateElements_0;
    SBox5Stage_mul2Context_delay_47_stateElements_1 <= SBox5Stage_mul2Context_delay_46_stateElements_1;
    SBox5Stage_mul2Context_delay_47_stateElements_2 <= SBox5Stage_mul2Context_delay_46_stateElements_2;
    SBox5Stage_mul2Context_delay_47_stateElements_3 <= SBox5Stage_mul2Context_delay_46_stateElements_3;
    SBox5Stage_mul2Context_delay_47_stateElements_4 <= SBox5Stage_mul2Context_delay_46_stateElements_4;
    SBox5Stage_mul2Context_delay_47_stateElements_5 <= SBox5Stage_mul2Context_delay_46_stateElements_5;
    SBox5Stage_mul2Context_delay_47_stateElements_6 <= SBox5Stage_mul2Context_delay_46_stateElements_6;
    SBox5Stage_mul2Context_delay_47_stateElements_7 <= SBox5Stage_mul2Context_delay_46_stateElements_7;
    SBox5Stage_mul2Context_delay_47_stateElements_8 <= SBox5Stage_mul2Context_delay_46_stateElements_8;
    SBox5Stage_mul2Context_delay_47_stateElements_9 <= SBox5Stage_mul2Context_delay_46_stateElements_9;
    SBox5Stage_mul2Context_delay_47_stateElements_10 <= SBox5Stage_mul2Context_delay_46_stateElements_10;
    SBox5Stage_mul2Context_delay_48_isFull <= SBox5Stage_mul2Context_delay_47_isFull;
    SBox5Stage_mul2Context_delay_48_fullRound <= SBox5Stage_mul2Context_delay_47_fullRound;
    SBox5Stage_mul2Context_delay_48_partialRound <= SBox5Stage_mul2Context_delay_47_partialRound;
    SBox5Stage_mul2Context_delay_48_stateIndex <= SBox5Stage_mul2Context_delay_47_stateIndex;
    SBox5Stage_mul2Context_delay_48_stateSize <= SBox5Stage_mul2Context_delay_47_stateSize;
    SBox5Stage_mul2Context_delay_48_stateID <= SBox5Stage_mul2Context_delay_47_stateID;
    SBox5Stage_mul2Context_delay_48_stateElements_0 <= SBox5Stage_mul2Context_delay_47_stateElements_0;
    SBox5Stage_mul2Context_delay_48_stateElements_1 <= SBox5Stage_mul2Context_delay_47_stateElements_1;
    SBox5Stage_mul2Context_delay_48_stateElements_2 <= SBox5Stage_mul2Context_delay_47_stateElements_2;
    SBox5Stage_mul2Context_delay_48_stateElements_3 <= SBox5Stage_mul2Context_delay_47_stateElements_3;
    SBox5Stage_mul2Context_delay_48_stateElements_4 <= SBox5Stage_mul2Context_delay_47_stateElements_4;
    SBox5Stage_mul2Context_delay_48_stateElements_5 <= SBox5Stage_mul2Context_delay_47_stateElements_5;
    SBox5Stage_mul2Context_delay_48_stateElements_6 <= SBox5Stage_mul2Context_delay_47_stateElements_6;
    SBox5Stage_mul2Context_delay_48_stateElements_7 <= SBox5Stage_mul2Context_delay_47_stateElements_7;
    SBox5Stage_mul2Context_delay_48_stateElements_8 <= SBox5Stage_mul2Context_delay_47_stateElements_8;
    SBox5Stage_mul2Context_delay_48_stateElements_9 <= SBox5Stage_mul2Context_delay_47_stateElements_9;
    SBox5Stage_mul2Context_delay_48_stateElements_10 <= SBox5Stage_mul2Context_delay_47_stateElements_10;
    SBox5Stage_tempContext2_isFull <= SBox5Stage_mul2Context_delay_48_isFull;
    SBox5Stage_tempContext2_fullRound <= SBox5Stage_mul2Context_delay_48_fullRound;
    SBox5Stage_tempContext2_partialRound <= SBox5Stage_mul2Context_delay_48_partialRound;
    SBox5Stage_tempContext2_stateIndex <= SBox5Stage_mul2Context_delay_48_stateIndex;
    SBox5Stage_tempContext2_stateSize <= SBox5Stage_mul2Context_delay_48_stateSize;
    SBox5Stage_tempContext2_stateID <= SBox5Stage_mul2Context_delay_48_stateID;
    SBox5Stage_tempContext2_stateElements_0 <= SBox5Stage_mul2Context_delay_48_stateElements_0;
    SBox5Stage_tempContext2_stateElements_1 <= SBox5Stage_mul2Context_delay_48_stateElements_1;
    SBox5Stage_tempContext2_stateElements_2 <= SBox5Stage_mul2Context_delay_48_stateElements_2;
    SBox5Stage_tempContext2_stateElements_3 <= SBox5Stage_mul2Context_delay_48_stateElements_3;
    SBox5Stage_tempContext2_stateElements_4 <= SBox5Stage_mul2Context_delay_48_stateElements_4;
    SBox5Stage_tempContext2_stateElements_5 <= SBox5Stage_mul2Context_delay_48_stateElements_5;
    SBox5Stage_tempContext2_stateElements_6 <= SBox5Stage_mul2Context_delay_48_stateElements_6;
    SBox5Stage_tempContext2_stateElements_7 <= SBox5Stage_mul2Context_delay_48_stateElements_7;
    SBox5Stage_tempContext2_stateElements_8 <= SBox5Stage_mul2Context_delay_48_stateElements_8;
    SBox5Stage_tempContext2_stateElements_9 <= SBox5Stage_mul2Context_delay_48_stateElements_9;
    SBox5Stage_tempContext2_stateElements_10 <= SBox5Stage_mul2Context_delay_48_stateElements_10;
    AddRoundConstantStage_adderContext_delay_1_isFull <= AddRoundConstantStage_adderContext_isFull;
    AddRoundConstantStage_adderContext_delay_1_fullRound <= AddRoundConstantStage_adderContext_fullRound;
    AddRoundConstantStage_adderContext_delay_1_partialRound <= AddRoundConstantStage_adderContext_partialRound;
    AddRoundConstantStage_adderContext_delay_1_stateIndex <= AddRoundConstantStage_adderContext_stateIndex;
    AddRoundConstantStage_adderContext_delay_1_stateSize <= AddRoundConstantStage_adderContext_stateSize;
    AddRoundConstantStage_adderContext_delay_1_stateID <= AddRoundConstantStage_adderContext_stateID;
    AddRoundConstantStage_adderContext_delay_1_stateElements_0 <= AddRoundConstantStage_adderContext_stateElements_0;
    AddRoundConstantStage_adderContext_delay_1_stateElements_1 <= AddRoundConstantStage_adderContext_stateElements_1;
    AddRoundConstantStage_adderContext_delay_1_stateElements_2 <= AddRoundConstantStage_adderContext_stateElements_2;
    AddRoundConstantStage_adderContext_delay_1_stateElements_3 <= AddRoundConstantStage_adderContext_stateElements_3;
    AddRoundConstantStage_adderContext_delay_1_stateElements_4 <= AddRoundConstantStage_adderContext_stateElements_4;
    AddRoundConstantStage_adderContext_delay_1_stateElements_5 <= AddRoundConstantStage_adderContext_stateElements_5;
    AddRoundConstantStage_adderContext_delay_1_stateElements_6 <= AddRoundConstantStage_adderContext_stateElements_6;
    AddRoundConstantStage_adderContext_delay_1_stateElements_7 <= AddRoundConstantStage_adderContext_stateElements_7;
    AddRoundConstantStage_adderContext_delay_1_stateElements_8 <= AddRoundConstantStage_adderContext_stateElements_8;
    AddRoundConstantStage_adderContext_delay_1_stateElements_9 <= AddRoundConstantStage_adderContext_stateElements_9;
    AddRoundConstantStage_adderContext_delay_1_stateElements_10 <= AddRoundConstantStage_adderContext_stateElements_10;
    AddRoundConstantStage_adderContext_delay_2_isFull <= AddRoundConstantStage_adderContext_delay_1_isFull;
    AddRoundConstantStage_adderContext_delay_2_fullRound <= AddRoundConstantStage_adderContext_delay_1_fullRound;
    AddRoundConstantStage_adderContext_delay_2_partialRound <= AddRoundConstantStage_adderContext_delay_1_partialRound;
    AddRoundConstantStage_adderContext_delay_2_stateIndex <= AddRoundConstantStage_adderContext_delay_1_stateIndex;
    AddRoundConstantStage_adderContext_delay_2_stateSize <= AddRoundConstantStage_adderContext_delay_1_stateSize;
    AddRoundConstantStage_adderContext_delay_2_stateID <= AddRoundConstantStage_adderContext_delay_1_stateID;
    AddRoundConstantStage_adderContext_delay_2_stateElements_0 <= AddRoundConstantStage_adderContext_delay_1_stateElements_0;
    AddRoundConstantStage_adderContext_delay_2_stateElements_1 <= AddRoundConstantStage_adderContext_delay_1_stateElements_1;
    AddRoundConstantStage_adderContext_delay_2_stateElements_2 <= AddRoundConstantStage_adderContext_delay_1_stateElements_2;
    AddRoundConstantStage_adderContext_delay_2_stateElements_3 <= AddRoundConstantStage_adderContext_delay_1_stateElements_3;
    AddRoundConstantStage_adderContext_delay_2_stateElements_4 <= AddRoundConstantStage_adderContext_delay_1_stateElements_4;
    AddRoundConstantStage_adderContext_delay_2_stateElements_5 <= AddRoundConstantStage_adderContext_delay_1_stateElements_5;
    AddRoundConstantStage_adderContext_delay_2_stateElements_6 <= AddRoundConstantStage_adderContext_delay_1_stateElements_6;
    AddRoundConstantStage_adderContext_delay_2_stateElements_7 <= AddRoundConstantStage_adderContext_delay_1_stateElements_7;
    AddRoundConstantStage_adderContext_delay_2_stateElements_8 <= AddRoundConstantStage_adderContext_delay_1_stateElements_8;
    AddRoundConstantStage_adderContext_delay_2_stateElements_9 <= AddRoundConstantStage_adderContext_delay_1_stateElements_9;
    AddRoundConstantStage_adderContext_delay_2_stateElements_10 <= AddRoundConstantStage_adderContext_delay_1_stateElements_10;
    AddRoundConstantStage_adderContext_delay_3_isFull <= AddRoundConstantStage_adderContext_delay_2_isFull;
    AddRoundConstantStage_adderContext_delay_3_fullRound <= AddRoundConstantStage_adderContext_delay_2_fullRound;
    AddRoundConstantStage_adderContext_delay_3_partialRound <= AddRoundConstantStage_adderContext_delay_2_partialRound;
    AddRoundConstantStage_adderContext_delay_3_stateIndex <= AddRoundConstantStage_adderContext_delay_2_stateIndex;
    AddRoundConstantStage_adderContext_delay_3_stateSize <= AddRoundConstantStage_adderContext_delay_2_stateSize;
    AddRoundConstantStage_adderContext_delay_3_stateID <= AddRoundConstantStage_adderContext_delay_2_stateID;
    AddRoundConstantStage_adderContext_delay_3_stateElements_0 <= AddRoundConstantStage_adderContext_delay_2_stateElements_0;
    AddRoundConstantStage_adderContext_delay_3_stateElements_1 <= AddRoundConstantStage_adderContext_delay_2_stateElements_1;
    AddRoundConstantStage_adderContext_delay_3_stateElements_2 <= AddRoundConstantStage_adderContext_delay_2_stateElements_2;
    AddRoundConstantStage_adderContext_delay_3_stateElements_3 <= AddRoundConstantStage_adderContext_delay_2_stateElements_3;
    AddRoundConstantStage_adderContext_delay_3_stateElements_4 <= AddRoundConstantStage_adderContext_delay_2_stateElements_4;
    AddRoundConstantStage_adderContext_delay_3_stateElements_5 <= AddRoundConstantStage_adderContext_delay_2_stateElements_5;
    AddRoundConstantStage_adderContext_delay_3_stateElements_6 <= AddRoundConstantStage_adderContext_delay_2_stateElements_6;
    AddRoundConstantStage_adderContext_delay_3_stateElements_7 <= AddRoundConstantStage_adderContext_delay_2_stateElements_7;
    AddRoundConstantStage_adderContext_delay_3_stateElements_8 <= AddRoundConstantStage_adderContext_delay_2_stateElements_8;
    AddRoundConstantStage_adderContext_delay_3_stateElements_9 <= AddRoundConstantStage_adderContext_delay_2_stateElements_9;
    AddRoundConstantStage_adderContext_delay_3_stateElements_10 <= AddRoundConstantStage_adderContext_delay_2_stateElements_10;
    AddRoundConstantStage_adderContext_delay_4_isFull <= AddRoundConstantStage_adderContext_delay_3_isFull;
    AddRoundConstantStage_adderContext_delay_4_fullRound <= AddRoundConstantStage_adderContext_delay_3_fullRound;
    AddRoundConstantStage_adderContext_delay_4_partialRound <= AddRoundConstantStage_adderContext_delay_3_partialRound;
    AddRoundConstantStage_adderContext_delay_4_stateIndex <= AddRoundConstantStage_adderContext_delay_3_stateIndex;
    AddRoundConstantStage_adderContext_delay_4_stateSize <= AddRoundConstantStage_adderContext_delay_3_stateSize;
    AddRoundConstantStage_adderContext_delay_4_stateID <= AddRoundConstantStage_adderContext_delay_3_stateID;
    AddRoundConstantStage_adderContext_delay_4_stateElements_0 <= AddRoundConstantStage_adderContext_delay_3_stateElements_0;
    AddRoundConstantStage_adderContext_delay_4_stateElements_1 <= AddRoundConstantStage_adderContext_delay_3_stateElements_1;
    AddRoundConstantStage_adderContext_delay_4_stateElements_2 <= AddRoundConstantStage_adderContext_delay_3_stateElements_2;
    AddRoundConstantStage_adderContext_delay_4_stateElements_3 <= AddRoundConstantStage_adderContext_delay_3_stateElements_3;
    AddRoundConstantStage_adderContext_delay_4_stateElements_4 <= AddRoundConstantStage_adderContext_delay_3_stateElements_4;
    AddRoundConstantStage_adderContext_delay_4_stateElements_5 <= AddRoundConstantStage_adderContext_delay_3_stateElements_5;
    AddRoundConstantStage_adderContext_delay_4_stateElements_6 <= AddRoundConstantStage_adderContext_delay_3_stateElements_6;
    AddRoundConstantStage_adderContext_delay_4_stateElements_7 <= AddRoundConstantStage_adderContext_delay_3_stateElements_7;
    AddRoundConstantStage_adderContext_delay_4_stateElements_8 <= AddRoundConstantStage_adderContext_delay_3_stateElements_8;
    AddRoundConstantStage_adderContext_delay_4_stateElements_9 <= AddRoundConstantStage_adderContext_delay_3_stateElements_9;
    AddRoundConstantStage_adderContext_delay_4_stateElements_10 <= AddRoundConstantStage_adderContext_delay_3_stateElements_10;
    AddRoundConstantStage_adderContext_delay_5_isFull <= AddRoundConstantStage_adderContext_delay_4_isFull;
    AddRoundConstantStage_adderContext_delay_5_fullRound <= AddRoundConstantStage_adderContext_delay_4_fullRound;
    AddRoundConstantStage_adderContext_delay_5_partialRound <= AddRoundConstantStage_adderContext_delay_4_partialRound;
    AddRoundConstantStage_adderContext_delay_5_stateIndex <= AddRoundConstantStage_adderContext_delay_4_stateIndex;
    AddRoundConstantStage_adderContext_delay_5_stateSize <= AddRoundConstantStage_adderContext_delay_4_stateSize;
    AddRoundConstantStage_adderContext_delay_5_stateID <= AddRoundConstantStage_adderContext_delay_4_stateID;
    AddRoundConstantStage_adderContext_delay_5_stateElements_0 <= AddRoundConstantStage_adderContext_delay_4_stateElements_0;
    AddRoundConstantStage_adderContext_delay_5_stateElements_1 <= AddRoundConstantStage_adderContext_delay_4_stateElements_1;
    AddRoundConstantStage_adderContext_delay_5_stateElements_2 <= AddRoundConstantStage_adderContext_delay_4_stateElements_2;
    AddRoundConstantStage_adderContext_delay_5_stateElements_3 <= AddRoundConstantStage_adderContext_delay_4_stateElements_3;
    AddRoundConstantStage_adderContext_delay_5_stateElements_4 <= AddRoundConstantStage_adderContext_delay_4_stateElements_4;
    AddRoundConstantStage_adderContext_delay_5_stateElements_5 <= AddRoundConstantStage_adderContext_delay_4_stateElements_5;
    AddRoundConstantStage_adderContext_delay_5_stateElements_6 <= AddRoundConstantStage_adderContext_delay_4_stateElements_6;
    AddRoundConstantStage_adderContext_delay_5_stateElements_7 <= AddRoundConstantStage_adderContext_delay_4_stateElements_7;
    AddRoundConstantStage_adderContext_delay_5_stateElements_8 <= AddRoundConstantStage_adderContext_delay_4_stateElements_8;
    AddRoundConstantStage_adderContext_delay_5_stateElements_9 <= AddRoundConstantStage_adderContext_delay_4_stateElements_9;
    AddRoundConstantStage_adderContext_delay_5_stateElements_10 <= AddRoundConstantStage_adderContext_delay_4_stateElements_10;
    AddRoundConstantStage_adderContext_delay_6_isFull <= AddRoundConstantStage_adderContext_delay_5_isFull;
    AddRoundConstantStage_adderContext_delay_6_fullRound <= AddRoundConstantStage_adderContext_delay_5_fullRound;
    AddRoundConstantStage_adderContext_delay_6_partialRound <= AddRoundConstantStage_adderContext_delay_5_partialRound;
    AddRoundConstantStage_adderContext_delay_6_stateIndex <= AddRoundConstantStage_adderContext_delay_5_stateIndex;
    AddRoundConstantStage_adderContext_delay_6_stateSize <= AddRoundConstantStage_adderContext_delay_5_stateSize;
    AddRoundConstantStage_adderContext_delay_6_stateID <= AddRoundConstantStage_adderContext_delay_5_stateID;
    AddRoundConstantStage_adderContext_delay_6_stateElements_0 <= AddRoundConstantStage_adderContext_delay_5_stateElements_0;
    AddRoundConstantStage_adderContext_delay_6_stateElements_1 <= AddRoundConstantStage_adderContext_delay_5_stateElements_1;
    AddRoundConstantStage_adderContext_delay_6_stateElements_2 <= AddRoundConstantStage_adderContext_delay_5_stateElements_2;
    AddRoundConstantStage_adderContext_delay_6_stateElements_3 <= AddRoundConstantStage_adderContext_delay_5_stateElements_3;
    AddRoundConstantStage_adderContext_delay_6_stateElements_4 <= AddRoundConstantStage_adderContext_delay_5_stateElements_4;
    AddRoundConstantStage_adderContext_delay_6_stateElements_5 <= AddRoundConstantStage_adderContext_delay_5_stateElements_5;
    AddRoundConstantStage_adderContext_delay_6_stateElements_6 <= AddRoundConstantStage_adderContext_delay_5_stateElements_6;
    AddRoundConstantStage_adderContext_delay_6_stateElements_7 <= AddRoundConstantStage_adderContext_delay_5_stateElements_7;
    AddRoundConstantStage_adderContext_delay_6_stateElements_8 <= AddRoundConstantStage_adderContext_delay_5_stateElements_8;
    AddRoundConstantStage_adderContext_delay_6_stateElements_9 <= AddRoundConstantStage_adderContext_delay_5_stateElements_9;
    AddRoundConstantStage_adderContext_delay_6_stateElements_10 <= AddRoundConstantStage_adderContext_delay_5_stateElements_10;
    AddRoundConstantStage_adderContext_delay_7_isFull <= AddRoundConstantStage_adderContext_delay_6_isFull;
    AddRoundConstantStage_adderContext_delay_7_fullRound <= AddRoundConstantStage_adderContext_delay_6_fullRound;
    AddRoundConstantStage_adderContext_delay_7_partialRound <= AddRoundConstantStage_adderContext_delay_6_partialRound;
    AddRoundConstantStage_adderContext_delay_7_stateIndex <= AddRoundConstantStage_adderContext_delay_6_stateIndex;
    AddRoundConstantStage_adderContext_delay_7_stateSize <= AddRoundConstantStage_adderContext_delay_6_stateSize;
    AddRoundConstantStage_adderContext_delay_7_stateID <= AddRoundConstantStage_adderContext_delay_6_stateID;
    AddRoundConstantStage_adderContext_delay_7_stateElements_0 <= AddRoundConstantStage_adderContext_delay_6_stateElements_0;
    AddRoundConstantStage_adderContext_delay_7_stateElements_1 <= AddRoundConstantStage_adderContext_delay_6_stateElements_1;
    AddRoundConstantStage_adderContext_delay_7_stateElements_2 <= AddRoundConstantStage_adderContext_delay_6_stateElements_2;
    AddRoundConstantStage_adderContext_delay_7_stateElements_3 <= AddRoundConstantStage_adderContext_delay_6_stateElements_3;
    AddRoundConstantStage_adderContext_delay_7_stateElements_4 <= AddRoundConstantStage_adderContext_delay_6_stateElements_4;
    AddRoundConstantStage_adderContext_delay_7_stateElements_5 <= AddRoundConstantStage_adderContext_delay_6_stateElements_5;
    AddRoundConstantStage_adderContext_delay_7_stateElements_6 <= AddRoundConstantStage_adderContext_delay_6_stateElements_6;
    AddRoundConstantStage_adderContext_delay_7_stateElements_7 <= AddRoundConstantStage_adderContext_delay_6_stateElements_7;
    AddRoundConstantStage_adderContext_delay_7_stateElements_8 <= AddRoundConstantStage_adderContext_delay_6_stateElements_8;
    AddRoundConstantStage_adderContext_delay_7_stateElements_9 <= AddRoundConstantStage_adderContext_delay_6_stateElements_9;
    AddRoundConstantStage_adderContext_delay_7_stateElements_10 <= AddRoundConstantStage_adderContext_delay_6_stateElements_10;
    AddRoundConstantStage_adderContext_delay_8_isFull <= AddRoundConstantStage_adderContext_delay_7_isFull;
    AddRoundConstantStage_adderContext_delay_8_fullRound <= AddRoundConstantStage_adderContext_delay_7_fullRound;
    AddRoundConstantStage_adderContext_delay_8_partialRound <= AddRoundConstantStage_adderContext_delay_7_partialRound;
    AddRoundConstantStage_adderContext_delay_8_stateIndex <= AddRoundConstantStage_adderContext_delay_7_stateIndex;
    AddRoundConstantStage_adderContext_delay_8_stateSize <= AddRoundConstantStage_adderContext_delay_7_stateSize;
    AddRoundConstantStage_adderContext_delay_8_stateID <= AddRoundConstantStage_adderContext_delay_7_stateID;
    AddRoundConstantStage_adderContext_delay_8_stateElements_0 <= AddRoundConstantStage_adderContext_delay_7_stateElements_0;
    AddRoundConstantStage_adderContext_delay_8_stateElements_1 <= AddRoundConstantStage_adderContext_delay_7_stateElements_1;
    AddRoundConstantStage_adderContext_delay_8_stateElements_2 <= AddRoundConstantStage_adderContext_delay_7_stateElements_2;
    AddRoundConstantStage_adderContext_delay_8_stateElements_3 <= AddRoundConstantStage_adderContext_delay_7_stateElements_3;
    AddRoundConstantStage_adderContext_delay_8_stateElements_4 <= AddRoundConstantStage_adderContext_delay_7_stateElements_4;
    AddRoundConstantStage_adderContext_delay_8_stateElements_5 <= AddRoundConstantStage_adderContext_delay_7_stateElements_5;
    AddRoundConstantStage_adderContext_delay_8_stateElements_6 <= AddRoundConstantStage_adderContext_delay_7_stateElements_6;
    AddRoundConstantStage_adderContext_delay_8_stateElements_7 <= AddRoundConstantStage_adderContext_delay_7_stateElements_7;
    AddRoundConstantStage_adderContext_delay_8_stateElements_8 <= AddRoundConstantStage_adderContext_delay_7_stateElements_8;
    AddRoundConstantStage_adderContext_delay_8_stateElements_9 <= AddRoundConstantStage_adderContext_delay_7_stateElements_9;
    AddRoundConstantStage_adderContext_delay_8_stateElements_10 <= AddRoundConstantStage_adderContext_delay_7_stateElements_10;
    AddRoundConstantStage_adderContext_delay_9_isFull <= AddRoundConstantStage_adderContext_delay_8_isFull;
    AddRoundConstantStage_adderContext_delay_9_fullRound <= AddRoundConstantStage_adderContext_delay_8_fullRound;
    AddRoundConstantStage_adderContext_delay_9_partialRound <= AddRoundConstantStage_adderContext_delay_8_partialRound;
    AddRoundConstantStage_adderContext_delay_9_stateIndex <= AddRoundConstantStage_adderContext_delay_8_stateIndex;
    AddRoundConstantStage_adderContext_delay_9_stateSize <= AddRoundConstantStage_adderContext_delay_8_stateSize;
    AddRoundConstantStage_adderContext_delay_9_stateID <= AddRoundConstantStage_adderContext_delay_8_stateID;
    AddRoundConstantStage_adderContext_delay_9_stateElements_0 <= AddRoundConstantStage_adderContext_delay_8_stateElements_0;
    AddRoundConstantStage_adderContext_delay_9_stateElements_1 <= AddRoundConstantStage_adderContext_delay_8_stateElements_1;
    AddRoundConstantStage_adderContext_delay_9_stateElements_2 <= AddRoundConstantStage_adderContext_delay_8_stateElements_2;
    AddRoundConstantStage_adderContext_delay_9_stateElements_3 <= AddRoundConstantStage_adderContext_delay_8_stateElements_3;
    AddRoundConstantStage_adderContext_delay_9_stateElements_4 <= AddRoundConstantStage_adderContext_delay_8_stateElements_4;
    AddRoundConstantStage_adderContext_delay_9_stateElements_5 <= AddRoundConstantStage_adderContext_delay_8_stateElements_5;
    AddRoundConstantStage_adderContext_delay_9_stateElements_6 <= AddRoundConstantStage_adderContext_delay_8_stateElements_6;
    AddRoundConstantStage_adderContext_delay_9_stateElements_7 <= AddRoundConstantStage_adderContext_delay_8_stateElements_7;
    AddRoundConstantStage_adderContext_delay_9_stateElements_8 <= AddRoundConstantStage_adderContext_delay_8_stateElements_8;
    AddRoundConstantStage_adderContext_delay_9_stateElements_9 <= AddRoundConstantStage_adderContext_delay_8_stateElements_9;
    AddRoundConstantStage_adderContext_delay_9_stateElements_10 <= AddRoundConstantStage_adderContext_delay_8_stateElements_10;
    AddRoundConstantStage_adderContext_delay_10_isFull <= AddRoundConstantStage_adderContext_delay_9_isFull;
    AddRoundConstantStage_adderContext_delay_10_fullRound <= AddRoundConstantStage_adderContext_delay_9_fullRound;
    AddRoundConstantStage_adderContext_delay_10_partialRound <= AddRoundConstantStage_adderContext_delay_9_partialRound;
    AddRoundConstantStage_adderContext_delay_10_stateIndex <= AddRoundConstantStage_adderContext_delay_9_stateIndex;
    AddRoundConstantStage_adderContext_delay_10_stateSize <= AddRoundConstantStage_adderContext_delay_9_stateSize;
    AddRoundConstantStage_adderContext_delay_10_stateID <= AddRoundConstantStage_adderContext_delay_9_stateID;
    AddRoundConstantStage_adderContext_delay_10_stateElements_0 <= AddRoundConstantStage_adderContext_delay_9_stateElements_0;
    AddRoundConstantStage_adderContext_delay_10_stateElements_1 <= AddRoundConstantStage_adderContext_delay_9_stateElements_1;
    AddRoundConstantStage_adderContext_delay_10_stateElements_2 <= AddRoundConstantStage_adderContext_delay_9_stateElements_2;
    AddRoundConstantStage_adderContext_delay_10_stateElements_3 <= AddRoundConstantStage_adderContext_delay_9_stateElements_3;
    AddRoundConstantStage_adderContext_delay_10_stateElements_4 <= AddRoundConstantStage_adderContext_delay_9_stateElements_4;
    AddRoundConstantStage_adderContext_delay_10_stateElements_5 <= AddRoundConstantStage_adderContext_delay_9_stateElements_5;
    AddRoundConstantStage_adderContext_delay_10_stateElements_6 <= AddRoundConstantStage_adderContext_delay_9_stateElements_6;
    AddRoundConstantStage_adderContext_delay_10_stateElements_7 <= AddRoundConstantStage_adderContext_delay_9_stateElements_7;
    AddRoundConstantStage_adderContext_delay_10_stateElements_8 <= AddRoundConstantStage_adderContext_delay_9_stateElements_8;
    AddRoundConstantStage_adderContext_delay_10_stateElements_9 <= AddRoundConstantStage_adderContext_delay_9_stateElements_9;
    AddRoundConstantStage_adderContext_delay_10_stateElements_10 <= AddRoundConstantStage_adderContext_delay_9_stateElements_10;
    AddRoundConstantStage_adderContext_delay_11_isFull <= AddRoundConstantStage_adderContext_delay_10_isFull;
    AddRoundConstantStage_adderContext_delay_11_fullRound <= AddRoundConstantStage_adderContext_delay_10_fullRound;
    AddRoundConstantStage_adderContext_delay_11_partialRound <= AddRoundConstantStage_adderContext_delay_10_partialRound;
    AddRoundConstantStage_adderContext_delay_11_stateIndex <= AddRoundConstantStage_adderContext_delay_10_stateIndex;
    AddRoundConstantStage_adderContext_delay_11_stateSize <= AddRoundConstantStage_adderContext_delay_10_stateSize;
    AddRoundConstantStage_adderContext_delay_11_stateID <= AddRoundConstantStage_adderContext_delay_10_stateID;
    AddRoundConstantStage_adderContext_delay_11_stateElements_0 <= AddRoundConstantStage_adderContext_delay_10_stateElements_0;
    AddRoundConstantStage_adderContext_delay_11_stateElements_1 <= AddRoundConstantStage_adderContext_delay_10_stateElements_1;
    AddRoundConstantStage_adderContext_delay_11_stateElements_2 <= AddRoundConstantStage_adderContext_delay_10_stateElements_2;
    AddRoundConstantStage_adderContext_delay_11_stateElements_3 <= AddRoundConstantStage_adderContext_delay_10_stateElements_3;
    AddRoundConstantStage_adderContext_delay_11_stateElements_4 <= AddRoundConstantStage_adderContext_delay_10_stateElements_4;
    AddRoundConstantStage_adderContext_delay_11_stateElements_5 <= AddRoundConstantStage_adderContext_delay_10_stateElements_5;
    AddRoundConstantStage_adderContext_delay_11_stateElements_6 <= AddRoundConstantStage_adderContext_delay_10_stateElements_6;
    AddRoundConstantStage_adderContext_delay_11_stateElements_7 <= AddRoundConstantStage_adderContext_delay_10_stateElements_7;
    AddRoundConstantStage_adderContext_delay_11_stateElements_8 <= AddRoundConstantStage_adderContext_delay_10_stateElements_8;
    AddRoundConstantStage_adderContext_delay_11_stateElements_9 <= AddRoundConstantStage_adderContext_delay_10_stateElements_9;
    AddRoundConstantStage_adderContext_delay_11_stateElements_10 <= AddRoundConstantStage_adderContext_delay_10_stateElements_10;
    AddRoundConstantStage_adderContext_delay_12_isFull <= AddRoundConstantStage_adderContext_delay_11_isFull;
    AddRoundConstantStage_adderContext_delay_12_fullRound <= AddRoundConstantStage_adderContext_delay_11_fullRound;
    AddRoundConstantStage_adderContext_delay_12_partialRound <= AddRoundConstantStage_adderContext_delay_11_partialRound;
    AddRoundConstantStage_adderContext_delay_12_stateIndex <= AddRoundConstantStage_adderContext_delay_11_stateIndex;
    AddRoundConstantStage_adderContext_delay_12_stateSize <= AddRoundConstantStage_adderContext_delay_11_stateSize;
    AddRoundConstantStage_adderContext_delay_12_stateID <= AddRoundConstantStage_adderContext_delay_11_stateID;
    AddRoundConstantStage_adderContext_delay_12_stateElements_0 <= AddRoundConstantStage_adderContext_delay_11_stateElements_0;
    AddRoundConstantStage_adderContext_delay_12_stateElements_1 <= AddRoundConstantStage_adderContext_delay_11_stateElements_1;
    AddRoundConstantStage_adderContext_delay_12_stateElements_2 <= AddRoundConstantStage_adderContext_delay_11_stateElements_2;
    AddRoundConstantStage_adderContext_delay_12_stateElements_3 <= AddRoundConstantStage_adderContext_delay_11_stateElements_3;
    AddRoundConstantStage_adderContext_delay_12_stateElements_4 <= AddRoundConstantStage_adderContext_delay_11_stateElements_4;
    AddRoundConstantStage_adderContext_delay_12_stateElements_5 <= AddRoundConstantStage_adderContext_delay_11_stateElements_5;
    AddRoundConstantStage_adderContext_delay_12_stateElements_6 <= AddRoundConstantStage_adderContext_delay_11_stateElements_6;
    AddRoundConstantStage_adderContext_delay_12_stateElements_7 <= AddRoundConstantStage_adderContext_delay_11_stateElements_7;
    AddRoundConstantStage_adderContext_delay_12_stateElements_8 <= AddRoundConstantStage_adderContext_delay_11_stateElements_8;
    AddRoundConstantStage_adderContext_delay_12_stateElements_9 <= AddRoundConstantStage_adderContext_delay_11_stateElements_9;
    AddRoundConstantStage_adderContext_delay_12_stateElements_10 <= AddRoundConstantStage_adderContext_delay_11_stateElements_10;
    AddRoundConstantStage_adderContext_delay_13_isFull <= AddRoundConstantStage_adderContext_delay_12_isFull;
    AddRoundConstantStage_adderContext_delay_13_fullRound <= AddRoundConstantStage_adderContext_delay_12_fullRound;
    AddRoundConstantStage_adderContext_delay_13_partialRound <= AddRoundConstantStage_adderContext_delay_12_partialRound;
    AddRoundConstantStage_adderContext_delay_13_stateIndex <= AddRoundConstantStage_adderContext_delay_12_stateIndex;
    AddRoundConstantStage_adderContext_delay_13_stateSize <= AddRoundConstantStage_adderContext_delay_12_stateSize;
    AddRoundConstantStage_adderContext_delay_13_stateID <= AddRoundConstantStage_adderContext_delay_12_stateID;
    AddRoundConstantStage_adderContext_delay_13_stateElements_0 <= AddRoundConstantStage_adderContext_delay_12_stateElements_0;
    AddRoundConstantStage_adderContext_delay_13_stateElements_1 <= AddRoundConstantStage_adderContext_delay_12_stateElements_1;
    AddRoundConstantStage_adderContext_delay_13_stateElements_2 <= AddRoundConstantStage_adderContext_delay_12_stateElements_2;
    AddRoundConstantStage_adderContext_delay_13_stateElements_3 <= AddRoundConstantStage_adderContext_delay_12_stateElements_3;
    AddRoundConstantStage_adderContext_delay_13_stateElements_4 <= AddRoundConstantStage_adderContext_delay_12_stateElements_4;
    AddRoundConstantStage_adderContext_delay_13_stateElements_5 <= AddRoundConstantStage_adderContext_delay_12_stateElements_5;
    AddRoundConstantStage_adderContext_delay_13_stateElements_6 <= AddRoundConstantStage_adderContext_delay_12_stateElements_6;
    AddRoundConstantStage_adderContext_delay_13_stateElements_7 <= AddRoundConstantStage_adderContext_delay_12_stateElements_7;
    AddRoundConstantStage_adderContext_delay_13_stateElements_8 <= AddRoundConstantStage_adderContext_delay_12_stateElements_8;
    AddRoundConstantStage_adderContext_delay_13_stateElements_9 <= AddRoundConstantStage_adderContext_delay_12_stateElements_9;
    AddRoundConstantStage_adderContext_delay_13_stateElements_10 <= AddRoundConstantStage_adderContext_delay_12_stateElements_10;
    AddRoundConstantStage_adderContext_delay_14_isFull <= AddRoundConstantStage_adderContext_delay_13_isFull;
    AddRoundConstantStage_adderContext_delay_14_fullRound <= AddRoundConstantStage_adderContext_delay_13_fullRound;
    AddRoundConstantStage_adderContext_delay_14_partialRound <= AddRoundConstantStage_adderContext_delay_13_partialRound;
    AddRoundConstantStage_adderContext_delay_14_stateIndex <= AddRoundConstantStage_adderContext_delay_13_stateIndex;
    AddRoundConstantStage_adderContext_delay_14_stateSize <= AddRoundConstantStage_adderContext_delay_13_stateSize;
    AddRoundConstantStage_adderContext_delay_14_stateID <= AddRoundConstantStage_adderContext_delay_13_stateID;
    AddRoundConstantStage_adderContext_delay_14_stateElements_0 <= AddRoundConstantStage_adderContext_delay_13_stateElements_0;
    AddRoundConstantStage_adderContext_delay_14_stateElements_1 <= AddRoundConstantStage_adderContext_delay_13_stateElements_1;
    AddRoundConstantStage_adderContext_delay_14_stateElements_2 <= AddRoundConstantStage_adderContext_delay_13_stateElements_2;
    AddRoundConstantStage_adderContext_delay_14_stateElements_3 <= AddRoundConstantStage_adderContext_delay_13_stateElements_3;
    AddRoundConstantStage_adderContext_delay_14_stateElements_4 <= AddRoundConstantStage_adderContext_delay_13_stateElements_4;
    AddRoundConstantStage_adderContext_delay_14_stateElements_5 <= AddRoundConstantStage_adderContext_delay_13_stateElements_5;
    AddRoundConstantStage_adderContext_delay_14_stateElements_6 <= AddRoundConstantStage_adderContext_delay_13_stateElements_6;
    AddRoundConstantStage_adderContext_delay_14_stateElements_7 <= AddRoundConstantStage_adderContext_delay_13_stateElements_7;
    AddRoundConstantStage_adderContext_delay_14_stateElements_8 <= AddRoundConstantStage_adderContext_delay_13_stateElements_8;
    AddRoundConstantStage_adderContext_delay_14_stateElements_9 <= AddRoundConstantStage_adderContext_delay_13_stateElements_9;
    AddRoundConstantStage_adderContext_delay_14_stateElements_10 <= AddRoundConstantStage_adderContext_delay_13_stateElements_10;
    AddRoundConstantStage_adderContext_delay_15_isFull <= AddRoundConstantStage_adderContext_delay_14_isFull;
    AddRoundConstantStage_adderContext_delay_15_fullRound <= AddRoundConstantStage_adderContext_delay_14_fullRound;
    AddRoundConstantStage_adderContext_delay_15_partialRound <= AddRoundConstantStage_adderContext_delay_14_partialRound;
    AddRoundConstantStage_adderContext_delay_15_stateIndex <= AddRoundConstantStage_adderContext_delay_14_stateIndex;
    AddRoundConstantStage_adderContext_delay_15_stateSize <= AddRoundConstantStage_adderContext_delay_14_stateSize;
    AddRoundConstantStage_adderContext_delay_15_stateID <= AddRoundConstantStage_adderContext_delay_14_stateID;
    AddRoundConstantStage_adderContext_delay_15_stateElements_0 <= AddRoundConstantStage_adderContext_delay_14_stateElements_0;
    AddRoundConstantStage_adderContext_delay_15_stateElements_1 <= AddRoundConstantStage_adderContext_delay_14_stateElements_1;
    AddRoundConstantStage_adderContext_delay_15_stateElements_2 <= AddRoundConstantStage_adderContext_delay_14_stateElements_2;
    AddRoundConstantStage_adderContext_delay_15_stateElements_3 <= AddRoundConstantStage_adderContext_delay_14_stateElements_3;
    AddRoundConstantStage_adderContext_delay_15_stateElements_4 <= AddRoundConstantStage_adderContext_delay_14_stateElements_4;
    AddRoundConstantStage_adderContext_delay_15_stateElements_5 <= AddRoundConstantStage_adderContext_delay_14_stateElements_5;
    AddRoundConstantStage_adderContext_delay_15_stateElements_6 <= AddRoundConstantStage_adderContext_delay_14_stateElements_6;
    AddRoundConstantStage_adderContext_delay_15_stateElements_7 <= AddRoundConstantStage_adderContext_delay_14_stateElements_7;
    AddRoundConstantStage_adderContext_delay_15_stateElements_8 <= AddRoundConstantStage_adderContext_delay_14_stateElements_8;
    AddRoundConstantStage_adderContext_delay_15_stateElements_9 <= AddRoundConstantStage_adderContext_delay_14_stateElements_9;
    AddRoundConstantStage_adderContext_delay_15_stateElements_10 <= AddRoundConstantStage_adderContext_delay_14_stateElements_10;
    AddRoundConstantStage_adderContext_delay_16_isFull <= AddRoundConstantStage_adderContext_delay_15_isFull;
    AddRoundConstantStage_adderContext_delay_16_fullRound <= AddRoundConstantStage_adderContext_delay_15_fullRound;
    AddRoundConstantStage_adderContext_delay_16_partialRound <= AddRoundConstantStage_adderContext_delay_15_partialRound;
    AddRoundConstantStage_adderContext_delay_16_stateIndex <= AddRoundConstantStage_adderContext_delay_15_stateIndex;
    AddRoundConstantStage_adderContext_delay_16_stateSize <= AddRoundConstantStage_adderContext_delay_15_stateSize;
    AddRoundConstantStage_adderContext_delay_16_stateID <= AddRoundConstantStage_adderContext_delay_15_stateID;
    AddRoundConstantStage_adderContext_delay_16_stateElements_0 <= AddRoundConstantStage_adderContext_delay_15_stateElements_0;
    AddRoundConstantStage_adderContext_delay_16_stateElements_1 <= AddRoundConstantStage_adderContext_delay_15_stateElements_1;
    AddRoundConstantStage_adderContext_delay_16_stateElements_2 <= AddRoundConstantStage_adderContext_delay_15_stateElements_2;
    AddRoundConstantStage_adderContext_delay_16_stateElements_3 <= AddRoundConstantStage_adderContext_delay_15_stateElements_3;
    AddRoundConstantStage_adderContext_delay_16_stateElements_4 <= AddRoundConstantStage_adderContext_delay_15_stateElements_4;
    AddRoundConstantStage_adderContext_delay_16_stateElements_5 <= AddRoundConstantStage_adderContext_delay_15_stateElements_5;
    AddRoundConstantStage_adderContext_delay_16_stateElements_6 <= AddRoundConstantStage_adderContext_delay_15_stateElements_6;
    AddRoundConstantStage_adderContext_delay_16_stateElements_7 <= AddRoundConstantStage_adderContext_delay_15_stateElements_7;
    AddRoundConstantStage_adderContext_delay_16_stateElements_8 <= AddRoundConstantStage_adderContext_delay_15_stateElements_8;
    AddRoundConstantStage_adderContext_delay_16_stateElements_9 <= AddRoundConstantStage_adderContext_delay_15_stateElements_9;
    AddRoundConstantStage_adderContext_delay_16_stateElements_10 <= AddRoundConstantStage_adderContext_delay_15_stateElements_10;
    AddRoundConstantStage_adderContext_delay_17_isFull <= AddRoundConstantStage_adderContext_delay_16_isFull;
    AddRoundConstantStage_adderContext_delay_17_fullRound <= AddRoundConstantStage_adderContext_delay_16_fullRound;
    AddRoundConstantStage_adderContext_delay_17_partialRound <= AddRoundConstantStage_adderContext_delay_16_partialRound;
    AddRoundConstantStage_adderContext_delay_17_stateIndex <= AddRoundConstantStage_adderContext_delay_16_stateIndex;
    AddRoundConstantStage_adderContext_delay_17_stateSize <= AddRoundConstantStage_adderContext_delay_16_stateSize;
    AddRoundConstantStage_adderContext_delay_17_stateID <= AddRoundConstantStage_adderContext_delay_16_stateID;
    AddRoundConstantStage_adderContext_delay_17_stateElements_0 <= AddRoundConstantStage_adderContext_delay_16_stateElements_0;
    AddRoundConstantStage_adderContext_delay_17_stateElements_1 <= AddRoundConstantStage_adderContext_delay_16_stateElements_1;
    AddRoundConstantStage_adderContext_delay_17_stateElements_2 <= AddRoundConstantStage_adderContext_delay_16_stateElements_2;
    AddRoundConstantStage_adderContext_delay_17_stateElements_3 <= AddRoundConstantStage_adderContext_delay_16_stateElements_3;
    AddRoundConstantStage_adderContext_delay_17_stateElements_4 <= AddRoundConstantStage_adderContext_delay_16_stateElements_4;
    AddRoundConstantStage_adderContext_delay_17_stateElements_5 <= AddRoundConstantStage_adderContext_delay_16_stateElements_5;
    AddRoundConstantStage_adderContext_delay_17_stateElements_6 <= AddRoundConstantStage_adderContext_delay_16_stateElements_6;
    AddRoundConstantStage_adderContext_delay_17_stateElements_7 <= AddRoundConstantStage_adderContext_delay_16_stateElements_7;
    AddRoundConstantStage_adderContext_delay_17_stateElements_8 <= AddRoundConstantStage_adderContext_delay_16_stateElements_8;
    AddRoundConstantStage_adderContext_delay_17_stateElements_9 <= AddRoundConstantStage_adderContext_delay_16_stateElements_9;
    AddRoundConstantStage_adderContext_delay_17_stateElements_10 <= AddRoundConstantStage_adderContext_delay_16_stateElements_10;
    AddRoundConstantStage_adderContext_delay_18_isFull <= AddRoundConstantStage_adderContext_delay_17_isFull;
    AddRoundConstantStage_adderContext_delay_18_fullRound <= AddRoundConstantStage_adderContext_delay_17_fullRound;
    AddRoundConstantStage_adderContext_delay_18_partialRound <= AddRoundConstantStage_adderContext_delay_17_partialRound;
    AddRoundConstantStage_adderContext_delay_18_stateIndex <= AddRoundConstantStage_adderContext_delay_17_stateIndex;
    AddRoundConstantStage_adderContext_delay_18_stateSize <= AddRoundConstantStage_adderContext_delay_17_stateSize;
    AddRoundConstantStage_adderContext_delay_18_stateID <= AddRoundConstantStage_adderContext_delay_17_stateID;
    AddRoundConstantStage_adderContext_delay_18_stateElements_0 <= AddRoundConstantStage_adderContext_delay_17_stateElements_0;
    AddRoundConstantStage_adderContext_delay_18_stateElements_1 <= AddRoundConstantStage_adderContext_delay_17_stateElements_1;
    AddRoundConstantStage_adderContext_delay_18_stateElements_2 <= AddRoundConstantStage_adderContext_delay_17_stateElements_2;
    AddRoundConstantStage_adderContext_delay_18_stateElements_3 <= AddRoundConstantStage_adderContext_delay_17_stateElements_3;
    AddRoundConstantStage_adderContext_delay_18_stateElements_4 <= AddRoundConstantStage_adderContext_delay_17_stateElements_4;
    AddRoundConstantStage_adderContext_delay_18_stateElements_5 <= AddRoundConstantStage_adderContext_delay_17_stateElements_5;
    AddRoundConstantStage_adderContext_delay_18_stateElements_6 <= AddRoundConstantStage_adderContext_delay_17_stateElements_6;
    AddRoundConstantStage_adderContext_delay_18_stateElements_7 <= AddRoundConstantStage_adderContext_delay_17_stateElements_7;
    AddRoundConstantStage_adderContext_delay_18_stateElements_8 <= AddRoundConstantStage_adderContext_delay_17_stateElements_8;
    AddRoundConstantStage_adderContext_delay_18_stateElements_9 <= AddRoundConstantStage_adderContext_delay_17_stateElements_9;
    AddRoundConstantStage_adderContext_delay_18_stateElements_10 <= AddRoundConstantStage_adderContext_delay_17_stateElements_10;
    AddRoundConstantStage_adderContext_delay_19_isFull <= AddRoundConstantStage_adderContext_delay_18_isFull;
    AddRoundConstantStage_adderContext_delay_19_fullRound <= AddRoundConstantStage_adderContext_delay_18_fullRound;
    AddRoundConstantStage_adderContext_delay_19_partialRound <= AddRoundConstantStage_adderContext_delay_18_partialRound;
    AddRoundConstantStage_adderContext_delay_19_stateIndex <= AddRoundConstantStage_adderContext_delay_18_stateIndex;
    AddRoundConstantStage_adderContext_delay_19_stateSize <= AddRoundConstantStage_adderContext_delay_18_stateSize;
    AddRoundConstantStage_adderContext_delay_19_stateID <= AddRoundConstantStage_adderContext_delay_18_stateID;
    AddRoundConstantStage_adderContext_delay_19_stateElements_0 <= AddRoundConstantStage_adderContext_delay_18_stateElements_0;
    AddRoundConstantStage_adderContext_delay_19_stateElements_1 <= AddRoundConstantStage_adderContext_delay_18_stateElements_1;
    AddRoundConstantStage_adderContext_delay_19_stateElements_2 <= AddRoundConstantStage_adderContext_delay_18_stateElements_2;
    AddRoundConstantStage_adderContext_delay_19_stateElements_3 <= AddRoundConstantStage_adderContext_delay_18_stateElements_3;
    AddRoundConstantStage_adderContext_delay_19_stateElements_4 <= AddRoundConstantStage_adderContext_delay_18_stateElements_4;
    AddRoundConstantStage_adderContext_delay_19_stateElements_5 <= AddRoundConstantStage_adderContext_delay_18_stateElements_5;
    AddRoundConstantStage_adderContext_delay_19_stateElements_6 <= AddRoundConstantStage_adderContext_delay_18_stateElements_6;
    AddRoundConstantStage_adderContext_delay_19_stateElements_7 <= AddRoundConstantStage_adderContext_delay_18_stateElements_7;
    AddRoundConstantStage_adderContext_delay_19_stateElements_8 <= AddRoundConstantStage_adderContext_delay_18_stateElements_8;
    AddRoundConstantStage_adderContext_delay_19_stateElements_9 <= AddRoundConstantStage_adderContext_delay_18_stateElements_9;
    AddRoundConstantStage_adderContext_delay_19_stateElements_10 <= AddRoundConstantStage_adderContext_delay_18_stateElements_10;
    AddRoundConstantStage_adderContext_delay_20_isFull <= AddRoundConstantStage_adderContext_delay_19_isFull;
    AddRoundConstantStage_adderContext_delay_20_fullRound <= AddRoundConstantStage_adderContext_delay_19_fullRound;
    AddRoundConstantStage_adderContext_delay_20_partialRound <= AddRoundConstantStage_adderContext_delay_19_partialRound;
    AddRoundConstantStage_adderContext_delay_20_stateIndex <= AddRoundConstantStage_adderContext_delay_19_stateIndex;
    AddRoundConstantStage_adderContext_delay_20_stateSize <= AddRoundConstantStage_adderContext_delay_19_stateSize;
    AddRoundConstantStage_adderContext_delay_20_stateID <= AddRoundConstantStage_adderContext_delay_19_stateID;
    AddRoundConstantStage_adderContext_delay_20_stateElements_0 <= AddRoundConstantStage_adderContext_delay_19_stateElements_0;
    AddRoundConstantStage_adderContext_delay_20_stateElements_1 <= AddRoundConstantStage_adderContext_delay_19_stateElements_1;
    AddRoundConstantStage_adderContext_delay_20_stateElements_2 <= AddRoundConstantStage_adderContext_delay_19_stateElements_2;
    AddRoundConstantStage_adderContext_delay_20_stateElements_3 <= AddRoundConstantStage_adderContext_delay_19_stateElements_3;
    AddRoundConstantStage_adderContext_delay_20_stateElements_4 <= AddRoundConstantStage_adderContext_delay_19_stateElements_4;
    AddRoundConstantStage_adderContext_delay_20_stateElements_5 <= AddRoundConstantStage_adderContext_delay_19_stateElements_5;
    AddRoundConstantStage_adderContext_delay_20_stateElements_6 <= AddRoundConstantStage_adderContext_delay_19_stateElements_6;
    AddRoundConstantStage_adderContext_delay_20_stateElements_7 <= AddRoundConstantStage_adderContext_delay_19_stateElements_7;
    AddRoundConstantStage_adderContext_delay_20_stateElements_8 <= AddRoundConstantStage_adderContext_delay_19_stateElements_8;
    AddRoundConstantStage_adderContext_delay_20_stateElements_9 <= AddRoundConstantStage_adderContext_delay_19_stateElements_9;
    AddRoundConstantStage_adderContext_delay_20_stateElements_10 <= AddRoundConstantStage_adderContext_delay_19_stateElements_10;
    AddRoundConstantStage_adderContext_delay_21_isFull <= AddRoundConstantStage_adderContext_delay_20_isFull;
    AddRoundConstantStage_adderContext_delay_21_fullRound <= AddRoundConstantStage_adderContext_delay_20_fullRound;
    AddRoundConstantStage_adderContext_delay_21_partialRound <= AddRoundConstantStage_adderContext_delay_20_partialRound;
    AddRoundConstantStage_adderContext_delay_21_stateIndex <= AddRoundConstantStage_adderContext_delay_20_stateIndex;
    AddRoundConstantStage_adderContext_delay_21_stateSize <= AddRoundConstantStage_adderContext_delay_20_stateSize;
    AddRoundConstantStage_adderContext_delay_21_stateID <= AddRoundConstantStage_adderContext_delay_20_stateID;
    AddRoundConstantStage_adderContext_delay_21_stateElements_0 <= AddRoundConstantStage_adderContext_delay_20_stateElements_0;
    AddRoundConstantStage_adderContext_delay_21_stateElements_1 <= AddRoundConstantStage_adderContext_delay_20_stateElements_1;
    AddRoundConstantStage_adderContext_delay_21_stateElements_2 <= AddRoundConstantStage_adderContext_delay_20_stateElements_2;
    AddRoundConstantStage_adderContext_delay_21_stateElements_3 <= AddRoundConstantStage_adderContext_delay_20_stateElements_3;
    AddRoundConstantStage_adderContext_delay_21_stateElements_4 <= AddRoundConstantStage_adderContext_delay_20_stateElements_4;
    AddRoundConstantStage_adderContext_delay_21_stateElements_5 <= AddRoundConstantStage_adderContext_delay_20_stateElements_5;
    AddRoundConstantStage_adderContext_delay_21_stateElements_6 <= AddRoundConstantStage_adderContext_delay_20_stateElements_6;
    AddRoundConstantStage_adderContext_delay_21_stateElements_7 <= AddRoundConstantStage_adderContext_delay_20_stateElements_7;
    AddRoundConstantStage_adderContext_delay_21_stateElements_8 <= AddRoundConstantStage_adderContext_delay_20_stateElements_8;
    AddRoundConstantStage_adderContext_delay_21_stateElements_9 <= AddRoundConstantStage_adderContext_delay_20_stateElements_9;
    AddRoundConstantStage_adderContext_delay_21_stateElements_10 <= AddRoundConstantStage_adderContext_delay_20_stateElements_10;
    AddRoundConstantStage_adderContext_delay_22_isFull <= AddRoundConstantStage_adderContext_delay_21_isFull;
    AddRoundConstantStage_adderContext_delay_22_fullRound <= AddRoundConstantStage_adderContext_delay_21_fullRound;
    AddRoundConstantStage_adderContext_delay_22_partialRound <= AddRoundConstantStage_adderContext_delay_21_partialRound;
    AddRoundConstantStage_adderContext_delay_22_stateIndex <= AddRoundConstantStage_adderContext_delay_21_stateIndex;
    AddRoundConstantStage_adderContext_delay_22_stateSize <= AddRoundConstantStage_adderContext_delay_21_stateSize;
    AddRoundConstantStage_adderContext_delay_22_stateID <= AddRoundConstantStage_adderContext_delay_21_stateID;
    AddRoundConstantStage_adderContext_delay_22_stateElements_0 <= AddRoundConstantStage_adderContext_delay_21_stateElements_0;
    AddRoundConstantStage_adderContext_delay_22_stateElements_1 <= AddRoundConstantStage_adderContext_delay_21_stateElements_1;
    AddRoundConstantStage_adderContext_delay_22_stateElements_2 <= AddRoundConstantStage_adderContext_delay_21_stateElements_2;
    AddRoundConstantStage_adderContext_delay_22_stateElements_3 <= AddRoundConstantStage_adderContext_delay_21_stateElements_3;
    AddRoundConstantStage_adderContext_delay_22_stateElements_4 <= AddRoundConstantStage_adderContext_delay_21_stateElements_4;
    AddRoundConstantStage_adderContext_delay_22_stateElements_5 <= AddRoundConstantStage_adderContext_delay_21_stateElements_5;
    AddRoundConstantStage_adderContext_delay_22_stateElements_6 <= AddRoundConstantStage_adderContext_delay_21_stateElements_6;
    AddRoundConstantStage_adderContext_delay_22_stateElements_7 <= AddRoundConstantStage_adderContext_delay_21_stateElements_7;
    AddRoundConstantStage_adderContext_delay_22_stateElements_8 <= AddRoundConstantStage_adderContext_delay_21_stateElements_8;
    AddRoundConstantStage_adderContext_delay_22_stateElements_9 <= AddRoundConstantStage_adderContext_delay_21_stateElements_9;
    AddRoundConstantStage_adderContext_delay_22_stateElements_10 <= AddRoundConstantStage_adderContext_delay_21_stateElements_10;
    AddRoundConstantStage_adderContext_delay_23_isFull <= AddRoundConstantStage_adderContext_delay_22_isFull;
    AddRoundConstantStage_adderContext_delay_23_fullRound <= AddRoundConstantStage_adderContext_delay_22_fullRound;
    AddRoundConstantStage_adderContext_delay_23_partialRound <= AddRoundConstantStage_adderContext_delay_22_partialRound;
    AddRoundConstantStage_adderContext_delay_23_stateIndex <= AddRoundConstantStage_adderContext_delay_22_stateIndex;
    AddRoundConstantStage_adderContext_delay_23_stateSize <= AddRoundConstantStage_adderContext_delay_22_stateSize;
    AddRoundConstantStage_adderContext_delay_23_stateID <= AddRoundConstantStage_adderContext_delay_22_stateID;
    AddRoundConstantStage_adderContext_delay_23_stateElements_0 <= AddRoundConstantStage_adderContext_delay_22_stateElements_0;
    AddRoundConstantStage_adderContext_delay_23_stateElements_1 <= AddRoundConstantStage_adderContext_delay_22_stateElements_1;
    AddRoundConstantStage_adderContext_delay_23_stateElements_2 <= AddRoundConstantStage_adderContext_delay_22_stateElements_2;
    AddRoundConstantStage_adderContext_delay_23_stateElements_3 <= AddRoundConstantStage_adderContext_delay_22_stateElements_3;
    AddRoundConstantStage_adderContext_delay_23_stateElements_4 <= AddRoundConstantStage_adderContext_delay_22_stateElements_4;
    AddRoundConstantStage_adderContext_delay_23_stateElements_5 <= AddRoundConstantStage_adderContext_delay_22_stateElements_5;
    AddRoundConstantStage_adderContext_delay_23_stateElements_6 <= AddRoundConstantStage_adderContext_delay_22_stateElements_6;
    AddRoundConstantStage_adderContext_delay_23_stateElements_7 <= AddRoundConstantStage_adderContext_delay_22_stateElements_7;
    AddRoundConstantStage_adderContext_delay_23_stateElements_8 <= AddRoundConstantStage_adderContext_delay_22_stateElements_8;
    AddRoundConstantStage_adderContext_delay_23_stateElements_9 <= AddRoundConstantStage_adderContext_delay_22_stateElements_9;
    AddRoundConstantStage_adderContext_delay_23_stateElements_10 <= AddRoundConstantStage_adderContext_delay_22_stateElements_10;
    AddRoundConstantStage_adderContext_delay_24_isFull <= AddRoundConstantStage_adderContext_delay_23_isFull;
    AddRoundConstantStage_adderContext_delay_24_fullRound <= AddRoundConstantStage_adderContext_delay_23_fullRound;
    AddRoundConstantStage_adderContext_delay_24_partialRound <= AddRoundConstantStage_adderContext_delay_23_partialRound;
    AddRoundConstantStage_adderContext_delay_24_stateIndex <= AddRoundConstantStage_adderContext_delay_23_stateIndex;
    AddRoundConstantStage_adderContext_delay_24_stateSize <= AddRoundConstantStage_adderContext_delay_23_stateSize;
    AddRoundConstantStage_adderContext_delay_24_stateID <= AddRoundConstantStage_adderContext_delay_23_stateID;
    AddRoundConstantStage_adderContext_delay_24_stateElements_0 <= AddRoundConstantStage_adderContext_delay_23_stateElements_0;
    AddRoundConstantStage_adderContext_delay_24_stateElements_1 <= AddRoundConstantStage_adderContext_delay_23_stateElements_1;
    AddRoundConstantStage_adderContext_delay_24_stateElements_2 <= AddRoundConstantStage_adderContext_delay_23_stateElements_2;
    AddRoundConstantStage_adderContext_delay_24_stateElements_3 <= AddRoundConstantStage_adderContext_delay_23_stateElements_3;
    AddRoundConstantStage_adderContext_delay_24_stateElements_4 <= AddRoundConstantStage_adderContext_delay_23_stateElements_4;
    AddRoundConstantStage_adderContext_delay_24_stateElements_5 <= AddRoundConstantStage_adderContext_delay_23_stateElements_5;
    AddRoundConstantStage_adderContext_delay_24_stateElements_6 <= AddRoundConstantStage_adderContext_delay_23_stateElements_6;
    AddRoundConstantStage_adderContext_delay_24_stateElements_7 <= AddRoundConstantStage_adderContext_delay_23_stateElements_7;
    AddRoundConstantStage_adderContext_delay_24_stateElements_8 <= AddRoundConstantStage_adderContext_delay_23_stateElements_8;
    AddRoundConstantStage_adderContext_delay_24_stateElements_9 <= AddRoundConstantStage_adderContext_delay_23_stateElements_9;
    AddRoundConstantStage_adderContext_delay_24_stateElements_10 <= AddRoundConstantStage_adderContext_delay_23_stateElements_10;
    AddRoundConstantStage_adderContext_delay_25_isFull <= AddRoundConstantStage_adderContext_delay_24_isFull;
    AddRoundConstantStage_adderContext_delay_25_fullRound <= AddRoundConstantStage_adderContext_delay_24_fullRound;
    AddRoundConstantStage_adderContext_delay_25_partialRound <= AddRoundConstantStage_adderContext_delay_24_partialRound;
    AddRoundConstantStage_adderContext_delay_25_stateIndex <= AddRoundConstantStage_adderContext_delay_24_stateIndex;
    AddRoundConstantStage_adderContext_delay_25_stateSize <= AddRoundConstantStage_adderContext_delay_24_stateSize;
    AddRoundConstantStage_adderContext_delay_25_stateID <= AddRoundConstantStage_adderContext_delay_24_stateID;
    AddRoundConstantStage_adderContext_delay_25_stateElements_0 <= AddRoundConstantStage_adderContext_delay_24_stateElements_0;
    AddRoundConstantStage_adderContext_delay_25_stateElements_1 <= AddRoundConstantStage_adderContext_delay_24_stateElements_1;
    AddRoundConstantStage_adderContext_delay_25_stateElements_2 <= AddRoundConstantStage_adderContext_delay_24_stateElements_2;
    AddRoundConstantStage_adderContext_delay_25_stateElements_3 <= AddRoundConstantStage_adderContext_delay_24_stateElements_3;
    AddRoundConstantStage_adderContext_delay_25_stateElements_4 <= AddRoundConstantStage_adderContext_delay_24_stateElements_4;
    AddRoundConstantStage_adderContext_delay_25_stateElements_5 <= AddRoundConstantStage_adderContext_delay_24_stateElements_5;
    AddRoundConstantStage_adderContext_delay_25_stateElements_6 <= AddRoundConstantStage_adderContext_delay_24_stateElements_6;
    AddRoundConstantStage_adderContext_delay_25_stateElements_7 <= AddRoundConstantStage_adderContext_delay_24_stateElements_7;
    AddRoundConstantStage_adderContext_delay_25_stateElements_8 <= AddRoundConstantStage_adderContext_delay_24_stateElements_8;
    AddRoundConstantStage_adderContext_delay_25_stateElements_9 <= AddRoundConstantStage_adderContext_delay_24_stateElements_9;
    AddRoundConstantStage_adderContext_delay_25_stateElements_10 <= AddRoundConstantStage_adderContext_delay_24_stateElements_10;
    AddRoundConstantStage_adderContext_delay_26_isFull <= AddRoundConstantStage_adderContext_delay_25_isFull;
    AddRoundConstantStage_adderContext_delay_26_fullRound <= AddRoundConstantStage_adderContext_delay_25_fullRound;
    AddRoundConstantStage_adderContext_delay_26_partialRound <= AddRoundConstantStage_adderContext_delay_25_partialRound;
    AddRoundConstantStage_adderContext_delay_26_stateIndex <= AddRoundConstantStage_adderContext_delay_25_stateIndex;
    AddRoundConstantStage_adderContext_delay_26_stateSize <= AddRoundConstantStage_adderContext_delay_25_stateSize;
    AddRoundConstantStage_adderContext_delay_26_stateID <= AddRoundConstantStage_adderContext_delay_25_stateID;
    AddRoundConstantStage_adderContext_delay_26_stateElements_0 <= AddRoundConstantStage_adderContext_delay_25_stateElements_0;
    AddRoundConstantStage_adderContext_delay_26_stateElements_1 <= AddRoundConstantStage_adderContext_delay_25_stateElements_1;
    AddRoundConstantStage_adderContext_delay_26_stateElements_2 <= AddRoundConstantStage_adderContext_delay_25_stateElements_2;
    AddRoundConstantStage_adderContext_delay_26_stateElements_3 <= AddRoundConstantStage_adderContext_delay_25_stateElements_3;
    AddRoundConstantStage_adderContext_delay_26_stateElements_4 <= AddRoundConstantStage_adderContext_delay_25_stateElements_4;
    AddRoundConstantStage_adderContext_delay_26_stateElements_5 <= AddRoundConstantStage_adderContext_delay_25_stateElements_5;
    AddRoundConstantStage_adderContext_delay_26_stateElements_6 <= AddRoundConstantStage_adderContext_delay_25_stateElements_6;
    AddRoundConstantStage_adderContext_delay_26_stateElements_7 <= AddRoundConstantStage_adderContext_delay_25_stateElements_7;
    AddRoundConstantStage_adderContext_delay_26_stateElements_8 <= AddRoundConstantStage_adderContext_delay_25_stateElements_8;
    AddRoundConstantStage_adderContext_delay_26_stateElements_9 <= AddRoundConstantStage_adderContext_delay_25_stateElements_9;
    AddRoundConstantStage_adderContext_delay_26_stateElements_10 <= AddRoundConstantStage_adderContext_delay_25_stateElements_10;
    AddRoundConstantStage_adderContext_delay_27_isFull <= AddRoundConstantStage_adderContext_delay_26_isFull;
    AddRoundConstantStage_adderContext_delay_27_fullRound <= AddRoundConstantStage_adderContext_delay_26_fullRound;
    AddRoundConstantStage_adderContext_delay_27_partialRound <= AddRoundConstantStage_adderContext_delay_26_partialRound;
    AddRoundConstantStage_adderContext_delay_27_stateIndex <= AddRoundConstantStage_adderContext_delay_26_stateIndex;
    AddRoundConstantStage_adderContext_delay_27_stateSize <= AddRoundConstantStage_adderContext_delay_26_stateSize;
    AddRoundConstantStage_adderContext_delay_27_stateID <= AddRoundConstantStage_adderContext_delay_26_stateID;
    AddRoundConstantStage_adderContext_delay_27_stateElements_0 <= AddRoundConstantStage_adderContext_delay_26_stateElements_0;
    AddRoundConstantStage_adderContext_delay_27_stateElements_1 <= AddRoundConstantStage_adderContext_delay_26_stateElements_1;
    AddRoundConstantStage_adderContext_delay_27_stateElements_2 <= AddRoundConstantStage_adderContext_delay_26_stateElements_2;
    AddRoundConstantStage_adderContext_delay_27_stateElements_3 <= AddRoundConstantStage_adderContext_delay_26_stateElements_3;
    AddRoundConstantStage_adderContext_delay_27_stateElements_4 <= AddRoundConstantStage_adderContext_delay_26_stateElements_4;
    AddRoundConstantStage_adderContext_delay_27_stateElements_5 <= AddRoundConstantStage_adderContext_delay_26_stateElements_5;
    AddRoundConstantStage_adderContext_delay_27_stateElements_6 <= AddRoundConstantStage_adderContext_delay_26_stateElements_6;
    AddRoundConstantStage_adderContext_delay_27_stateElements_7 <= AddRoundConstantStage_adderContext_delay_26_stateElements_7;
    AddRoundConstantStage_adderContext_delay_27_stateElements_8 <= AddRoundConstantStage_adderContext_delay_26_stateElements_8;
    AddRoundConstantStage_adderContext_delay_27_stateElements_9 <= AddRoundConstantStage_adderContext_delay_26_stateElements_9;
    AddRoundConstantStage_adderContext_delay_27_stateElements_10 <= AddRoundConstantStage_adderContext_delay_26_stateElements_10;
    AddRoundConstantStage_adderContext_delay_28_isFull <= AddRoundConstantStage_adderContext_delay_27_isFull;
    AddRoundConstantStage_adderContext_delay_28_fullRound <= AddRoundConstantStage_adderContext_delay_27_fullRound;
    AddRoundConstantStage_adderContext_delay_28_partialRound <= AddRoundConstantStage_adderContext_delay_27_partialRound;
    AddRoundConstantStage_adderContext_delay_28_stateIndex <= AddRoundConstantStage_adderContext_delay_27_stateIndex;
    AddRoundConstantStage_adderContext_delay_28_stateSize <= AddRoundConstantStage_adderContext_delay_27_stateSize;
    AddRoundConstantStage_adderContext_delay_28_stateID <= AddRoundConstantStage_adderContext_delay_27_stateID;
    AddRoundConstantStage_adderContext_delay_28_stateElements_0 <= AddRoundConstantStage_adderContext_delay_27_stateElements_0;
    AddRoundConstantStage_adderContext_delay_28_stateElements_1 <= AddRoundConstantStage_adderContext_delay_27_stateElements_1;
    AddRoundConstantStage_adderContext_delay_28_stateElements_2 <= AddRoundConstantStage_adderContext_delay_27_stateElements_2;
    AddRoundConstantStage_adderContext_delay_28_stateElements_3 <= AddRoundConstantStage_adderContext_delay_27_stateElements_3;
    AddRoundConstantStage_adderContext_delay_28_stateElements_4 <= AddRoundConstantStage_adderContext_delay_27_stateElements_4;
    AddRoundConstantStage_adderContext_delay_28_stateElements_5 <= AddRoundConstantStage_adderContext_delay_27_stateElements_5;
    AddRoundConstantStage_adderContext_delay_28_stateElements_6 <= AddRoundConstantStage_adderContext_delay_27_stateElements_6;
    AddRoundConstantStage_adderContext_delay_28_stateElements_7 <= AddRoundConstantStage_adderContext_delay_27_stateElements_7;
    AddRoundConstantStage_adderContext_delay_28_stateElements_8 <= AddRoundConstantStage_adderContext_delay_27_stateElements_8;
    AddRoundConstantStage_adderContext_delay_28_stateElements_9 <= AddRoundConstantStage_adderContext_delay_27_stateElements_9;
    AddRoundConstantStage_adderContext_delay_28_stateElements_10 <= AddRoundConstantStage_adderContext_delay_27_stateElements_10;
    AddRoundConstantStage_adderContext_delay_29_isFull <= AddRoundConstantStage_adderContext_delay_28_isFull;
    AddRoundConstantStage_adderContext_delay_29_fullRound <= AddRoundConstantStage_adderContext_delay_28_fullRound;
    AddRoundConstantStage_adderContext_delay_29_partialRound <= AddRoundConstantStage_adderContext_delay_28_partialRound;
    AddRoundConstantStage_adderContext_delay_29_stateIndex <= AddRoundConstantStage_adderContext_delay_28_stateIndex;
    AddRoundConstantStage_adderContext_delay_29_stateSize <= AddRoundConstantStage_adderContext_delay_28_stateSize;
    AddRoundConstantStage_adderContext_delay_29_stateID <= AddRoundConstantStage_adderContext_delay_28_stateID;
    AddRoundConstantStage_adderContext_delay_29_stateElements_0 <= AddRoundConstantStage_adderContext_delay_28_stateElements_0;
    AddRoundConstantStage_adderContext_delay_29_stateElements_1 <= AddRoundConstantStage_adderContext_delay_28_stateElements_1;
    AddRoundConstantStage_adderContext_delay_29_stateElements_2 <= AddRoundConstantStage_adderContext_delay_28_stateElements_2;
    AddRoundConstantStage_adderContext_delay_29_stateElements_3 <= AddRoundConstantStage_adderContext_delay_28_stateElements_3;
    AddRoundConstantStage_adderContext_delay_29_stateElements_4 <= AddRoundConstantStage_adderContext_delay_28_stateElements_4;
    AddRoundConstantStage_adderContext_delay_29_stateElements_5 <= AddRoundConstantStage_adderContext_delay_28_stateElements_5;
    AddRoundConstantStage_adderContext_delay_29_stateElements_6 <= AddRoundConstantStage_adderContext_delay_28_stateElements_6;
    AddRoundConstantStage_adderContext_delay_29_stateElements_7 <= AddRoundConstantStage_adderContext_delay_28_stateElements_7;
    AddRoundConstantStage_adderContext_delay_29_stateElements_8 <= AddRoundConstantStage_adderContext_delay_28_stateElements_8;
    AddRoundConstantStage_adderContext_delay_29_stateElements_9 <= AddRoundConstantStage_adderContext_delay_28_stateElements_9;
    AddRoundConstantStage_adderContext_delay_29_stateElements_10 <= AddRoundConstantStage_adderContext_delay_28_stateElements_10;
    AddRoundConstantStage_adderContext_delay_30_isFull <= AddRoundConstantStage_adderContext_delay_29_isFull;
    AddRoundConstantStage_adderContext_delay_30_fullRound <= AddRoundConstantStage_adderContext_delay_29_fullRound;
    AddRoundConstantStage_adderContext_delay_30_partialRound <= AddRoundConstantStage_adderContext_delay_29_partialRound;
    AddRoundConstantStage_adderContext_delay_30_stateIndex <= AddRoundConstantStage_adderContext_delay_29_stateIndex;
    AddRoundConstantStage_adderContext_delay_30_stateSize <= AddRoundConstantStage_adderContext_delay_29_stateSize;
    AddRoundConstantStage_adderContext_delay_30_stateID <= AddRoundConstantStage_adderContext_delay_29_stateID;
    AddRoundConstantStage_adderContext_delay_30_stateElements_0 <= AddRoundConstantStage_adderContext_delay_29_stateElements_0;
    AddRoundConstantStage_adderContext_delay_30_stateElements_1 <= AddRoundConstantStage_adderContext_delay_29_stateElements_1;
    AddRoundConstantStage_adderContext_delay_30_stateElements_2 <= AddRoundConstantStage_adderContext_delay_29_stateElements_2;
    AddRoundConstantStage_adderContext_delay_30_stateElements_3 <= AddRoundConstantStage_adderContext_delay_29_stateElements_3;
    AddRoundConstantStage_adderContext_delay_30_stateElements_4 <= AddRoundConstantStage_adderContext_delay_29_stateElements_4;
    AddRoundConstantStage_adderContext_delay_30_stateElements_5 <= AddRoundConstantStage_adderContext_delay_29_stateElements_5;
    AddRoundConstantStage_adderContext_delay_30_stateElements_6 <= AddRoundConstantStage_adderContext_delay_29_stateElements_6;
    AddRoundConstantStage_adderContext_delay_30_stateElements_7 <= AddRoundConstantStage_adderContext_delay_29_stateElements_7;
    AddRoundConstantStage_adderContext_delay_30_stateElements_8 <= AddRoundConstantStage_adderContext_delay_29_stateElements_8;
    AddRoundConstantStage_adderContext_delay_30_stateElements_9 <= AddRoundConstantStage_adderContext_delay_29_stateElements_9;
    AddRoundConstantStage_adderContext_delay_30_stateElements_10 <= AddRoundConstantStage_adderContext_delay_29_stateElements_10;
    AddRoundConstantStage_adderContext_delay_31_isFull <= AddRoundConstantStage_adderContext_delay_30_isFull;
    AddRoundConstantStage_adderContext_delay_31_fullRound <= AddRoundConstantStage_adderContext_delay_30_fullRound;
    AddRoundConstantStage_adderContext_delay_31_partialRound <= AddRoundConstantStage_adderContext_delay_30_partialRound;
    AddRoundConstantStage_adderContext_delay_31_stateIndex <= AddRoundConstantStage_adderContext_delay_30_stateIndex;
    AddRoundConstantStage_adderContext_delay_31_stateSize <= AddRoundConstantStage_adderContext_delay_30_stateSize;
    AddRoundConstantStage_adderContext_delay_31_stateID <= AddRoundConstantStage_adderContext_delay_30_stateID;
    AddRoundConstantStage_adderContext_delay_31_stateElements_0 <= AddRoundConstantStage_adderContext_delay_30_stateElements_0;
    AddRoundConstantStage_adderContext_delay_31_stateElements_1 <= AddRoundConstantStage_adderContext_delay_30_stateElements_1;
    AddRoundConstantStage_adderContext_delay_31_stateElements_2 <= AddRoundConstantStage_adderContext_delay_30_stateElements_2;
    AddRoundConstantStage_adderContext_delay_31_stateElements_3 <= AddRoundConstantStage_adderContext_delay_30_stateElements_3;
    AddRoundConstantStage_adderContext_delay_31_stateElements_4 <= AddRoundConstantStage_adderContext_delay_30_stateElements_4;
    AddRoundConstantStage_adderContext_delay_31_stateElements_5 <= AddRoundConstantStage_adderContext_delay_30_stateElements_5;
    AddRoundConstantStage_adderContext_delay_31_stateElements_6 <= AddRoundConstantStage_adderContext_delay_30_stateElements_6;
    AddRoundConstantStage_adderContext_delay_31_stateElements_7 <= AddRoundConstantStage_adderContext_delay_30_stateElements_7;
    AddRoundConstantStage_adderContext_delay_31_stateElements_8 <= AddRoundConstantStage_adderContext_delay_30_stateElements_8;
    AddRoundConstantStage_adderContext_delay_31_stateElements_9 <= AddRoundConstantStage_adderContext_delay_30_stateElements_9;
    AddRoundConstantStage_adderContext_delay_31_stateElements_10 <= AddRoundConstantStage_adderContext_delay_30_stateElements_10;
    AddRoundConstantStage_adderContext_delay_32_isFull <= AddRoundConstantStage_adderContext_delay_31_isFull;
    AddRoundConstantStage_adderContext_delay_32_fullRound <= AddRoundConstantStage_adderContext_delay_31_fullRound;
    AddRoundConstantStage_adderContext_delay_32_partialRound <= AddRoundConstantStage_adderContext_delay_31_partialRound;
    AddRoundConstantStage_adderContext_delay_32_stateIndex <= AddRoundConstantStage_adderContext_delay_31_stateIndex;
    AddRoundConstantStage_adderContext_delay_32_stateSize <= AddRoundConstantStage_adderContext_delay_31_stateSize;
    AddRoundConstantStage_adderContext_delay_32_stateID <= AddRoundConstantStage_adderContext_delay_31_stateID;
    AddRoundConstantStage_adderContext_delay_32_stateElements_0 <= AddRoundConstantStage_adderContext_delay_31_stateElements_0;
    AddRoundConstantStage_adderContext_delay_32_stateElements_1 <= AddRoundConstantStage_adderContext_delay_31_stateElements_1;
    AddRoundConstantStage_adderContext_delay_32_stateElements_2 <= AddRoundConstantStage_adderContext_delay_31_stateElements_2;
    AddRoundConstantStage_adderContext_delay_32_stateElements_3 <= AddRoundConstantStage_adderContext_delay_31_stateElements_3;
    AddRoundConstantStage_adderContext_delay_32_stateElements_4 <= AddRoundConstantStage_adderContext_delay_31_stateElements_4;
    AddRoundConstantStage_adderContext_delay_32_stateElements_5 <= AddRoundConstantStage_adderContext_delay_31_stateElements_5;
    AddRoundConstantStage_adderContext_delay_32_stateElements_6 <= AddRoundConstantStage_adderContext_delay_31_stateElements_6;
    AddRoundConstantStage_adderContext_delay_32_stateElements_7 <= AddRoundConstantStage_adderContext_delay_31_stateElements_7;
    AddRoundConstantStage_adderContext_delay_32_stateElements_8 <= AddRoundConstantStage_adderContext_delay_31_stateElements_8;
    AddRoundConstantStage_adderContext_delay_32_stateElements_9 <= AddRoundConstantStage_adderContext_delay_31_stateElements_9;
    AddRoundConstantStage_adderContext_delay_32_stateElements_10 <= AddRoundConstantStage_adderContext_delay_31_stateElements_10;
    AddRoundConstantStage_adderContextDelayed_isFull <= AddRoundConstantStage_adderContext_delay_32_isFull;
    AddRoundConstantStage_adderContextDelayed_fullRound <= AddRoundConstantStage_adderContext_delay_32_fullRound;
    AddRoundConstantStage_adderContextDelayed_partialRound <= AddRoundConstantStage_adderContext_delay_32_partialRound;
    AddRoundConstantStage_adderContextDelayed_stateIndex <= AddRoundConstantStage_adderContext_delay_32_stateIndex;
    AddRoundConstantStage_adderContextDelayed_stateSize <= AddRoundConstantStage_adderContext_delay_32_stateSize;
    AddRoundConstantStage_adderContextDelayed_stateID <= AddRoundConstantStage_adderContext_delay_32_stateID;
    AddRoundConstantStage_adderContextDelayed_stateElements_0 <= AddRoundConstantStage_adderContext_delay_32_stateElements_0;
    AddRoundConstantStage_adderContextDelayed_stateElements_1 <= AddRoundConstantStage_adderContext_delay_32_stateElements_1;
    AddRoundConstantStage_adderContextDelayed_stateElements_2 <= AddRoundConstantStage_adderContext_delay_32_stateElements_2;
    AddRoundConstantStage_adderContextDelayed_stateElements_3 <= AddRoundConstantStage_adderContext_delay_32_stateElements_3;
    AddRoundConstantStage_adderContextDelayed_stateElements_4 <= AddRoundConstantStage_adderContext_delay_32_stateElements_4;
    AddRoundConstantStage_adderContextDelayed_stateElements_5 <= AddRoundConstantStage_adderContext_delay_32_stateElements_5;
    AddRoundConstantStage_adderContextDelayed_stateElements_6 <= AddRoundConstantStage_adderContext_delay_32_stateElements_6;
    AddRoundConstantStage_adderContextDelayed_stateElements_7 <= AddRoundConstantStage_adderContext_delay_32_stateElements_7;
    AddRoundConstantStage_adderContextDelayed_stateElements_8 <= AddRoundConstantStage_adderContext_delay_32_stateElements_8;
    AddRoundConstantStage_adderContextDelayed_stateElements_9 <= AddRoundConstantStage_adderContext_delay_32_stateElements_9;
    AddRoundConstantStage_adderContextDelayed_stateElements_10 <= AddRoundConstantStage_adderContext_delay_32_stateElements_10;
    AddRoundConstantStage_output_regNext_payload_isFull <= AddRoundConstantStage_output_payload_isFull;
    AddRoundConstantStage_output_regNext_payload_fullRound <= AddRoundConstantStage_output_payload_fullRound;
    AddRoundConstantStage_output_regNext_payload_partialRound <= AddRoundConstantStage_output_payload_partialRound;
    AddRoundConstantStage_output_regNext_payload_stateIndex <= AddRoundConstantStage_output_payload_stateIndex;
    AddRoundConstantStage_output_regNext_payload_stateSize <= AddRoundConstantStage_output_payload_stateSize;
    AddRoundConstantStage_output_regNext_payload_stateID <= AddRoundConstantStage_output_payload_stateID;
    AddRoundConstantStage_output_regNext_payload_stateElements_0 <= AddRoundConstantStage_output_payload_stateElements_0;
    AddRoundConstantStage_output_regNext_payload_stateElements_1 <= AddRoundConstantStage_output_payload_stateElements_1;
    AddRoundConstantStage_output_regNext_payload_stateElements_2 <= AddRoundConstantStage_output_payload_stateElements_2;
    AddRoundConstantStage_output_regNext_payload_stateElements_3 <= AddRoundConstantStage_output_payload_stateElements_3;
    AddRoundConstantStage_output_regNext_payload_stateElements_4 <= AddRoundConstantStage_output_payload_stateElements_4;
    AddRoundConstantStage_output_regNext_payload_stateElements_5 <= AddRoundConstantStage_output_payload_stateElements_5;
    AddRoundConstantStage_output_regNext_payload_stateElements_6 <= AddRoundConstantStage_output_payload_stateElements_6;
    AddRoundConstantStage_output_regNext_payload_stateElements_7 <= AddRoundConstantStage_output_payload_stateElements_7;
    AddRoundConstantStage_output_regNext_payload_stateElements_8 <= AddRoundConstantStage_output_payload_stateElements_8;
    AddRoundConstantStage_output_regNext_payload_stateElements_9 <= AddRoundConstantStage_output_payload_stateElements_9;
    AddRoundConstantStage_output_regNext_payload_stateElements_10 <= AddRoundConstantStage_output_payload_stateElements_10;
    AddRoundConstantStage_output_regNext_payload_stateElement <= AddRoundConstantStage_output_payload_stateElement;
  end

  always @(posedge clk) begin
    if(!resetn) begin
      AddRoundConstantStage_output_regNext_valid <= 1'b0;
    end else begin
      AddRoundConstantStage_output_regNext_valid <= AddRoundConstantStage_output_valid;
    end
  end


endmodule

module ModularAdderFlow_1 (
  input               io_input_valid,
  input      [254:0]  io_input_payload_op1,
  input      [254:0]  io_input_payload_op2,
  output              io_output_valid,
  output     [254:0]  io_output_payload_res,
  input               clk,
  input               resetn
);

  wire                adderIPFlow_4_io_output_valid;
  wire       [255:0]  adderIPFlow_4_io_output_payload_res;
  wire                adderIPFlow_5_io_output_valid;
  wire       [255:0]  adderIPFlow_5_io_output_payload_res;
  wire       [255:0]  _zz__zz_io_output_payload_res;
  wire                adderInput2_valid;
  wire       [254:0]  adderInput2_payload_op1;
  wire       [254:0]  adderInput2_payload_op2;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_1;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_2;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_3;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_4;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_5;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_6;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_7;
  reg        [255:0]  res1Delayed;
  reg                 _zz_io_output_valid;
  reg        [254:0]  _zz_io_output_payload_res;

  assign _zz__zz_io_output_payload_res = ((adderIPFlow_5_io_output_payload_res[255] || res1Delayed[255]) ? adderIPFlow_5_io_output_payload_res : res1Delayed);
  AdderIPFlow_2 adderIPFlow_4 (
    .io_input_valid           (io_input_valid                              ), //i
    .io_input_payload_op1     (io_input_payload_op1[254:0]                 ), //i
    .io_input_payload_op2     (io_input_payload_op2[254:0]                 ), //i
    .io_output_valid          (adderIPFlow_4_io_output_valid               ), //o
    .io_output_payload_res    (adderIPFlow_4_io_output_payload_res[255:0]  ), //o
    .clk                      (clk                                         ), //i
    .resetn                   (resetn                                      )  //i
  );
  AdderIPFlow_2 adderIPFlow_5 (
    .io_input_valid           (adderInput2_valid                           ), //i
    .io_input_payload_op1     (adderInput2_payload_op1[254:0]              ), //i
    .io_input_payload_op2     (adderInput2_payload_op2[254:0]              ), //i
    .io_output_valid          (adderIPFlow_5_io_output_valid               ), //o
    .io_output_payload_res    (adderIPFlow_5_io_output_payload_res[255:0]  ), //o
    .clk                      (clk                                         ), //i
    .resetn                   (resetn                                      )  //i
  );
  assign adderInput2_valid = adderIPFlow_4_io_output_valid;
  assign adderInput2_payload_op1 = adderIPFlow_4_io_output_payload_res[254:0];
  assign adderInput2_payload_op2 = 255'h0c1258acd66282b7ccc627f7f65e27faac425bfd0001a40100000000ffffffff;
  assign io_output_valid = _zz_io_output_valid;
  assign io_output_payload_res = _zz_io_output_payload_res;
  always @(posedge clk) begin
    adderIPFlow_4_io_output_payload_res_delay_1 <= adderIPFlow_4_io_output_payload_res;
    adderIPFlow_4_io_output_payload_res_delay_2 <= adderIPFlow_4_io_output_payload_res_delay_1;
    adderIPFlow_4_io_output_payload_res_delay_3 <= adderIPFlow_4_io_output_payload_res_delay_2;
    adderIPFlow_4_io_output_payload_res_delay_4 <= adderIPFlow_4_io_output_payload_res_delay_3;
    adderIPFlow_4_io_output_payload_res_delay_5 <= adderIPFlow_4_io_output_payload_res_delay_4;
    adderIPFlow_4_io_output_payload_res_delay_6 <= adderIPFlow_4_io_output_payload_res_delay_5;
    adderIPFlow_4_io_output_payload_res_delay_7 <= adderIPFlow_4_io_output_payload_res_delay_6;
    res1Delayed <= adderIPFlow_4_io_output_payload_res_delay_7;
    _zz_io_output_payload_res <= _zz__zz_io_output_payload_res[254:0];
  end

  always @(posedge clk) begin
    if(!resetn) begin
      _zz_io_output_valid <= 1'b0;
    end else begin
      _zz_io_output_valid <= adderIPFlow_5_io_output_valid;
    end
  end


endmodule

module PreRoundConstantMem (
  input      [3:0]    io_stateSize,
  input      [3:0]    io_stateIndex,
  output     [254:0]  io_preConstant
);

  wire       [254:0]  _zz_memInst_0_port0;
  wire       [254:0]  _zz_memInst_1_port0;
  wire       [254:0]  _zz_memInst_2_port0;
  wire       [254:0]  _zz_memInst_3_port0;
  wire       [1:0]    _zz_memInst_0_port;
  wire       [1:0]    _zz_memOutput_0_1;
  wire       [2:0]    _zz_memInst_1_port;
  wire       [2:0]    _zz_memOutput_1_1;
  reg        [254:0]  _zz_io_preConstant_2;
  wire       [1:0]    _zz_io_preConstant_3;
  wire       [253:0]  initialContent_0_0;
  wire       [254:0]  initialContent_0_1;
  wire       [254:0]  initialContent_0_2;
  wire       [253:0]  initialContent_1_0;
  wire       [254:0]  initialContent_1_1;
  wire       [253:0]  initialContent_1_2;
  wire       [254:0]  initialContent_1_3;
  wire       [254:0]  initialContent_1_4;
  wire       [254:0]  initialContent_2_0;
  wire       [254:0]  initialContent_2_1;
  wire       [254:0]  initialContent_2_2;
  wire       [254:0]  initialContent_2_3;
  wire       [254:0]  initialContent_2_4;
  wire       [252:0]  initialContent_2_5;
  wire       [252:0]  initialContent_2_6;
  wire       [252:0]  initialContent_2_7;
  wire       [254:0]  initialContent_2_8;
  wire       [252:0]  initialContent_3_0;
  wire       [252:0]  initialContent_3_1;
  wire       [250:0]  initialContent_3_2;
  wire       [254:0]  initialContent_3_3;
  wire       [252:0]  initialContent_3_4;
  wire       [254:0]  initialContent_3_5;
  wire       [254:0]  initialContent_3_6;
  wire       [252:0]  initialContent_3_7;
  wire       [254:0]  initialContent_3_8;
  wire       [254:0]  initialContent_3_9;
  wire       [254:0]  initialContent_3_10;
  wire       [254:0]  initialContent_3_11;
  wire       [3:0]    _zz_memOutput_0;
  wire       [254:0]  memOutput_0;
  wire       [3:0]    _zz_memOutput_1;
  wire       [254:0]  memOutput_1;
  wire       [3:0]    _zz_memOutput_2;
  wire       [254:0]  memOutput_2;
  wire       [3:0]    _zz_memOutput_3;
  wire       [254:0]  memOutput_3;
  wire                select_0;
  wire                select_1;
  wire                select_2;
  wire                select_3;
  wire                _zz_io_preConstant;
  wire                _zz_io_preConstant_1;
  (* ram_style = "distributed" *) reg [254:0] memInst_0 [0:2];
  (* ram_style = "distributed" *) reg [254:0] memInst_1 [0:4];
  (* ram_style = "distributed" *) reg [254:0] memInst_2 [0:8];
  (* ram_style = "distributed" *) reg [254:0] memInst_3 [0:11];

  assign _zz_memOutput_0_1 = _zz_memOutput_0[1:0];
  assign _zz_memOutput_1_1 = _zz_memOutput_1[2:0];
  assign _zz_io_preConstant_3 = {_zz_io_preConstant_1,_zz_io_preConstant};
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_preRoundConstantMem_1_memInst_0.bin",memInst_0);
  end
  assign _zz_memInst_0_port0 = memInst_0[_zz_memOutput_0_1];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_preRoundConstantMem_1_memInst_1.bin",memInst_1);
  end
  assign _zz_memInst_1_port0 = memInst_1[_zz_memOutput_1_1];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_preRoundConstantMem_1_memInst_2.bin",memInst_2);
  end
  assign _zz_memInst_2_port0 = memInst_2[_zz_memOutput_2];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_preRoundConstantMem_1_memInst_3.bin",memInst_3);
  end
  assign _zz_memInst_3_port0 = memInst_3[_zz_memOutput_3];
  always @(*) begin
    case(_zz_io_preConstant_3)
      2'b00 : _zz_io_preConstant_2 = memOutput_0;
      2'b01 : _zz_io_preConstant_2 = memOutput_1;
      2'b10 : _zz_io_preConstant_2 = memOutput_2;
      default : _zz_io_preConstant_2 = memOutput_3;
    endcase
  end

  assign initialContent_0_0 = 254'h2a175464246e8941586440d29d17a3e801c1bdf20d09026b23e366d1c822c12d;
  assign initialContent_0_1 = 255'h600fd1b8363956cbdbfb4087da06af8ec28b6be869a2cf82dd35fb45585c6aed;
  assign initialContent_0_2 = 255'h69212d4e6495f3683deb63f13fe00e4249df84165dccb57f3fa379d7e2b8bfbe;
  assign initialContent_1_0 = 254'h33ff809e7dbdebbf8f644337a0008dcf305605b2cb53223d3d0a4729368cfb9f;
  assign initialContent_1_1 = 255'h4998feed41b4cddf2572ea256be885d0503170b7205090679e52ce58a4182072;
  assign initialContent_1_2 = 254'h27ae16683e3a7acc2302dadf7a5fa9c5034410574ac64bd6578b2978864d447c;
  assign initialContent_1_3 = 255'h5ec0e948c78bc2c24fbe333d330cfb35307db01f23092d8c6d3a7acd0bbd8dd7;
  assign initialContent_1_4 = 255'h73b33c1d097fe58c0b7c1572fafa5f3067d901cf30252eee2cb4d18b3637e7e5;
  assign initialContent_2_0 = 255'h61164ad53d961f8c5d71b17b8762cfe5b80a09c3770458818eb749221c5777b2;
  assign initialContent_2_1 = 255'h629457753f89131cd47ba9d8cd6946fe4d9710737560c27a773d3406a8f372e5;
  assign initialContent_2_2 = 255'h7107e746a7f5d03edf182e037acdc21dc049822362518bf52fcfc516572100c6;
  assign initialContent_2_3 = 255'h6d682d57c2f77a87982f101aa874cc41716286f9625d3d92a968983a5ef53811;
  assign initialContent_2_4 = 255'h5af7e3d8f26afd924b8d17a25ff21fe5e1d792d5f295095fb676e1da058ed62f;
  assign initialContent_2_5 = 253'h1df39ecbc80f8cd77fe8ecebd38a68bd8e96c48fda8e055c41b143e41b03fa28;
  assign initialContent_2_6 = 253'h130c8a1cdc46a1feaf252450edd7afc1810f5fe59bc15438855be06daacb38ca;
  assign initialContent_2_7 = 253'h1caed2dbef24448b570ba85bacd8d8a59674e1b0da119872e2a4a3fb359dcf90;
  assign initialContent_2_8 = 255'h5d2a5445b34a8c40f1642337f13047a2767d87551c943519380312717f01c615;
  assign initialContent_3_0 = 253'h17fa0c9a759f5b22f592e9170b46d35bec219c80c7f1f34d70bd48a2f2f6061f;
  assign initialContent_3_1 = 253'h1e380507358adb0dd4c8ff7007bd1f1f7fdf2350c0a4989b04f0d4cf72dc5c77;
  assign initialContent_3_2 = 251'h55baa6a9addd6703ae3a88059aeaf8176f3453533910eee7002dc13c81bfb07;
  assign initialContent_3_3 = 255'h59afa6e185c556f0c46834f185695aef105089c669bcebe48ffe7e848165e138;
  assign initialContent_3_4 = 253'h18e3e88a35ed841034d08f4c86633376a5404c484cf7e63bc4690dc8f2a12121;
  assign initialContent_3_5 = 255'h50f9329aad27d133c367c805dd6c5829ec24a9bd6d7a3cd9e7c46b528078d4d7;
  assign initialContent_3_6 = 255'h69a4eef12806819f181f6ba6aefe9cbe9c663618e7e8ba4c5a96cdeb798f7579;
  assign initialContent_3_7 = 253'h168c18dde57a2e4654bb324ccb241209c79ceb9b63830f21741b569b35071986;
  assign initialContent_3_8 = 255'h49f8d58a75a960d871dfd1ba40e985c10e39911645f5d35fadbffe3695ebab04;
  assign initialContent_3_9 = 255'h6163c52a1a4a5b5a4aad9cce14d6ffe6695d01abb6db317b877af0af830e804c;
  assign initialContent_3_10 = 255'h591b0c6bed72f4e6fdff7700591f2435b85c0361c6b226e2774779cdb0fc6d2e;
  assign initialContent_3_11 = 255'h586d4eacccd4167cf1538c8690df076bd88d48a64ea86aaecd6cda86c44450e0;
  assign _zz_memOutput_0 = io_stateIndex;
  assign memOutput_0 = _zz_memInst_0_port0;
  assign _zz_memOutput_1 = io_stateIndex;
  assign memOutput_1 = _zz_memInst_1_port0;
  assign _zz_memOutput_2 = io_stateIndex;
  assign memOutput_2 = _zz_memInst_2_port0;
  assign _zz_memOutput_3 = io_stateIndex;
  assign memOutput_3 = _zz_memInst_3_port0;
  assign select_0 = (io_stateSize == 4'b0011);
  assign select_1 = (io_stateSize == 4'b0101);
  assign select_2 = (io_stateSize == 4'b1001);
  assign select_3 = (io_stateSize == 4'b1100);
  assign _zz_io_preConstant = (select_1 || select_3);
  assign _zz_io_preConstant_1 = (select_2 || select_3);
  assign io_preConstant = _zz_io_preConstant_2;

endmodule

module PoseidonSerializer (
  input               io_input_valid,
  output reg          io_input_ready,
  input               io_input_payload_isFull,
  input      [2:0]    io_input_payload_fullRound,
  input      [5:0]    io_input_payload_partialRound,
  input      [3:0]    io_input_payload_stateSize,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElements_0,
  input      [254:0]  io_input_payload_stateElements_1,
  input      [254:0]  io_input_payload_stateElements_2,
  input      [254:0]  io_input_payload_stateElements_3,
  input      [254:0]  io_input_payload_stateElements_4,
  input      [254:0]  io_input_payload_stateElements_5,
  input      [254:0]  io_input_payload_stateElements_6,
  input      [254:0]  io_input_payload_stateElements_7,
  input      [254:0]  io_input_payload_stateElements_8,
  input      [254:0]  io_input_payload_stateElements_9,
  input      [254:0]  io_input_payload_stateElements_10,
  input      [254:0]  io_input_payload_stateElements_11,
  output reg          io_output_valid,
  input               io_output_ready,
  output              io_output_payload_isFull,
  output     [2:0]    io_output_payload_fullRound,
  output     [5:0]    io_output_payload_partialRound,
  output     [3:0]    io_output_payload_stateIndex,
  output     [3:0]    io_output_payload_stateSize,
  output     [7:0]    io_output_payload_stateID,
  output reg [254:0]  io_output_payload_stateElements_0,
  output reg [254:0]  io_output_payload_stateElements_1,
  output reg [254:0]  io_output_payload_stateElements_2,
  output reg [254:0]  io_output_payload_stateElements_3,
  output reg [254:0]  io_output_payload_stateElements_4,
  output reg [254:0]  io_output_payload_stateElements_5,
  output reg [254:0]  io_output_payload_stateElements_6,
  output reg [254:0]  io_output_payload_stateElements_7,
  output reg [254:0]  io_output_payload_stateElements_8,
  output reg [254:0]  io_output_payload_stateElements_9,
  output reg [254:0]  io_output_payload_stateElements_10,
  output reg [254:0]  io_output_payload_stateElement,
  input               clk,
  input               resetn
);
  localparam fsm_enumDef_BOOT = 3'd0;
  localparam fsm_enumDef_IDLE = 3'd1;
  localparam fsm_enumDef_FULL = 3'd2;
  localparam fsm_enumDef_PARTIAL = 3'd3;
  localparam fsm_enumDef_LAST = 3'd4;

  reg        [254:0]  _zz_io_output_payload_stateElement;
  wire       [3:0]    _zz_when_PoseidonSerializer_l73;
  reg                 buffer_isFull;
  reg        [2:0]    buffer_fullRound;
  reg        [5:0]    buffer_partialRound;
  reg        [3:0]    buffer_stateSize;
  reg        [7:0]    buffer_stateID;
  reg        [254:0]  buffer_stateElements_0;
  reg        [254:0]  buffer_stateElements_1;
  reg        [254:0]  buffer_stateElements_2;
  reg        [254:0]  buffer_stateElements_3;
  reg        [254:0]  buffer_stateElements_4;
  reg        [254:0]  buffer_stateElements_5;
  reg        [254:0]  buffer_stateElements_6;
  reg        [254:0]  buffer_stateElements_7;
  reg        [254:0]  buffer_stateElements_8;
  reg        [254:0]  buffer_stateElements_9;
  reg        [254:0]  buffer_stateElements_10;
  reg        [254:0]  buffer_stateElements_11;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg        [3:0]    fsm_counter;
  reg        [2:0]    fsm_stateReg;
  reg        [2:0]    fsm_stateNext;
  wire                io_input_fire;
  wire                when_PoseidonSerializer_l59;
  wire                io_output_fire;
  wire                when_PoseidonSerializer_l73;
  wire                io_output_fire_1;
  wire                when_PoseidonSerializer_l92;
  wire                io_output_fire_2;
  wire                io_input_fire_1;
  wire                when_PoseidonSerializer_l106;
  wire                when_StateMachine_l222;
  `ifndef SYNTHESIS
  reg [55:0] fsm_stateReg_string;
  reg [55:0] fsm_stateNext_string;
  `endif


  assign _zz_when_PoseidonSerializer_l73 = (buffer_stateSize - 4'b0010);
  always @(*) begin
    case(fsm_counter)
      4'b0000 : _zz_io_output_payload_stateElement = buffer_stateElements_0;
      4'b0001 : _zz_io_output_payload_stateElement = buffer_stateElements_1;
      4'b0010 : _zz_io_output_payload_stateElement = buffer_stateElements_2;
      4'b0011 : _zz_io_output_payload_stateElement = buffer_stateElements_3;
      4'b0100 : _zz_io_output_payload_stateElement = buffer_stateElements_4;
      4'b0101 : _zz_io_output_payload_stateElement = buffer_stateElements_5;
      4'b0110 : _zz_io_output_payload_stateElement = buffer_stateElements_6;
      4'b0111 : _zz_io_output_payload_stateElement = buffer_stateElements_7;
      4'b1000 : _zz_io_output_payload_stateElement = buffer_stateElements_8;
      4'b1001 : _zz_io_output_payload_stateElement = buffer_stateElements_9;
      4'b1010 : _zz_io_output_payload_stateElement = buffer_stateElements_10;
      default : _zz_io_output_payload_stateElement = buffer_stateElements_11;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_BOOT : fsm_stateReg_string = "BOOT   ";
      fsm_enumDef_IDLE : fsm_stateReg_string = "IDLE   ";
      fsm_enumDef_FULL : fsm_stateReg_string = "FULL   ";
      fsm_enumDef_PARTIAL : fsm_stateReg_string = "PARTIAL";
      fsm_enumDef_LAST : fsm_stateReg_string = "LAST   ";
      default : fsm_stateReg_string = "???????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_BOOT : fsm_stateNext_string = "BOOT   ";
      fsm_enumDef_IDLE : fsm_stateNext_string = "IDLE   ";
      fsm_enumDef_FULL : fsm_stateNext_string = "FULL   ";
      fsm_enumDef_PARTIAL : fsm_stateNext_string = "PARTIAL";
      fsm_enumDef_LAST : fsm_stateNext_string = "LAST   ";
      default : fsm_stateNext_string = "???????";
    endcase
  end
  `endif

  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
      end
      fsm_enumDef_LAST : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    io_input_ready = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
        io_input_ready = 1'b1;
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
      end
      fsm_enumDef_LAST : begin
        if(io_output_fire_2) begin
          io_input_ready = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_valid = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
        io_output_valid = 1'b1;
      end
      fsm_enumDef_PARTIAL : begin
        io_output_valid = 1'b1;
      end
      fsm_enumDef_LAST : begin
        io_output_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign io_output_payload_isFull = buffer_isFull;
  assign io_output_payload_fullRound = buffer_fullRound;
  assign io_output_payload_partialRound = buffer_partialRound;
  assign io_output_payload_stateIndex = fsm_counter;
  assign io_output_payload_stateSize = buffer_stateSize;
  assign io_output_payload_stateID = buffer_stateID;
  always @(*) begin
    io_output_payload_stateElement = _zz_io_output_payload_stateElement;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElement = buffer_stateElements_0;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_0 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_0 = buffer_stateElements_1;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_0 = buffer_stateElements_1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_1 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_1 = buffer_stateElements_2;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_1 = buffer_stateElements_2;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_2 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_2 = buffer_stateElements_3;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_2 = buffer_stateElements_3;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_3 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_3 = buffer_stateElements_4;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_3 = buffer_stateElements_4;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_4 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_4 = buffer_stateElements_5;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_4 = buffer_stateElements_5;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_5 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_5 = buffer_stateElements_6;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_5 = buffer_stateElements_6;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_6 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_6 = buffer_stateElements_7;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_6 = buffer_stateElements_7;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_7 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_7 = buffer_stateElements_8;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_7 = buffer_stateElements_8;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_8 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_8 = buffer_stateElements_9;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_8 = buffer_stateElements_9;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_9 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_9 = buffer_stateElements_10;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_9 = buffer_stateElements_10;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_10 = 255'h0;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
      end
      fsm_enumDef_FULL : begin
      end
      fsm_enumDef_PARTIAL : begin
        io_output_payload_stateElements_10 = buffer_stateElements_11;
      end
      fsm_enumDef_LAST : begin
        if(when_PoseidonSerializer_l92) begin
          io_output_payload_stateElements_10 = buffer_stateElements_11;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_IDLE : begin
        if(io_input_fire) begin
          if(io_input_payload_isFull) begin
            fsm_stateNext = fsm_enumDef_FULL;
          end else begin
            if(when_PoseidonSerializer_l59) begin
              fsm_stateNext = fsm_enumDef_LAST;
            end else begin
              fsm_stateNext = fsm_enumDef_PARTIAL;
            end
          end
        end
      end
      fsm_enumDef_FULL : begin
        if(io_output_fire) begin
          if(when_PoseidonSerializer_l73) begin
            fsm_stateNext = fsm_enumDef_LAST;
          end
        end
      end
      fsm_enumDef_PARTIAL : begin
        if(io_output_fire_1) begin
          fsm_stateNext = fsm_enumDef_LAST;
        end
      end
      fsm_enumDef_LAST : begin
        if(io_output_fire_2) begin
          if(io_input_fire_1) begin
            if(io_input_payload_isFull) begin
              fsm_stateNext = fsm_enumDef_FULL;
            end else begin
              if(when_PoseidonSerializer_l106) begin
                fsm_stateNext = fsm_enumDef_PARTIAL;
              end
            end
          end else begin
            fsm_stateNext = fsm_enumDef_IDLE;
          end
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_IDLE;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_BOOT;
    end
  end

  assign io_input_fire = (io_input_valid && io_input_ready);
  assign when_PoseidonSerializer_l59 = (io_input_payload_stateSize < 4'b1001);
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign when_PoseidonSerializer_l73 = (fsm_counter == _zz_when_PoseidonSerializer_l73);
  assign io_output_fire_1 = (io_output_valid && io_output_ready);
  assign when_PoseidonSerializer_l92 = (! buffer_isFull);
  assign io_output_fire_2 = (io_output_valid && io_output_ready);
  assign io_input_fire_1 = (io_input_valid && io_input_ready);
  assign when_PoseidonSerializer_l106 = (4'b0101 < io_input_payload_stateSize);
  assign when_StateMachine_l222 = ((fsm_stateReg == fsm_enumDef_LAST) && (! (fsm_stateNext == fsm_enumDef_LAST)));
  always @(posedge clk) begin
    if(!resetn) begin
      buffer_isFull <= 1'b0;
      buffer_fullRound <= 3'b000;
      buffer_partialRound <= 6'h0;
      buffer_stateSize <= 4'b0000;
      buffer_stateID <= 8'h0;
      buffer_stateElements_0 <= 255'h0;
      buffer_stateElements_1 <= 255'h0;
      buffer_stateElements_2 <= 255'h0;
      buffer_stateElements_3 <= 255'h0;
      buffer_stateElements_4 <= 255'h0;
      buffer_stateElements_5 <= 255'h0;
      buffer_stateElements_6 <= 255'h0;
      buffer_stateElements_7 <= 255'h0;
      buffer_stateElements_8 <= 255'h0;
      buffer_stateElements_9 <= 255'h0;
      buffer_stateElements_10 <= 255'h0;
      buffer_stateElements_11 <= 255'h0;
      fsm_counter <= 4'b0000;
      fsm_stateReg <= fsm_enumDef_BOOT;
    end else begin
      fsm_stateReg <= fsm_stateNext;
      case(fsm_stateReg)
        fsm_enumDef_IDLE : begin
          if(io_input_fire) begin
            buffer_isFull <= io_input_payload_isFull;
            buffer_fullRound <= io_input_payload_fullRound;
            buffer_partialRound <= io_input_payload_partialRound;
            buffer_stateSize <= io_input_payload_stateSize;
            buffer_stateID <= io_input_payload_stateID;
            buffer_stateElements_0 <= io_input_payload_stateElements_0;
            buffer_stateElements_1 <= io_input_payload_stateElements_1;
            buffer_stateElements_2 <= io_input_payload_stateElements_2;
            buffer_stateElements_3 <= io_input_payload_stateElements_3;
            buffer_stateElements_4 <= io_input_payload_stateElements_4;
            buffer_stateElements_5 <= io_input_payload_stateElements_5;
            buffer_stateElements_6 <= io_input_payload_stateElements_6;
            buffer_stateElements_7 <= io_input_payload_stateElements_7;
            buffer_stateElements_8 <= io_input_payload_stateElements_8;
            buffer_stateElements_9 <= io_input_payload_stateElements_9;
            buffer_stateElements_10 <= io_input_payload_stateElements_10;
            buffer_stateElements_11 <= io_input_payload_stateElements_11;
          end
        end
        fsm_enumDef_FULL : begin
          if(io_output_fire) begin
            fsm_counter <= (fsm_counter + 4'b0001);
          end
        end
        fsm_enumDef_PARTIAL : begin
          if(io_output_fire_1) begin
            fsm_counter <= (fsm_counter + 4'b0001);
          end
        end
        fsm_enumDef_LAST : begin
          if(io_output_fire_2) begin
            if(io_input_fire_1) begin
              buffer_isFull <= io_input_payload_isFull;
              buffer_fullRound <= io_input_payload_fullRound;
              buffer_partialRound <= io_input_payload_partialRound;
              buffer_stateSize <= io_input_payload_stateSize;
              buffer_stateID <= io_input_payload_stateID;
              buffer_stateElements_0 <= io_input_payload_stateElements_0;
              buffer_stateElements_1 <= io_input_payload_stateElements_1;
              buffer_stateElements_2 <= io_input_payload_stateElements_2;
              buffer_stateElements_3 <= io_input_payload_stateElements_3;
              buffer_stateElements_4 <= io_input_payload_stateElements_4;
              buffer_stateElements_5 <= io_input_payload_stateElements_5;
              buffer_stateElements_6 <= io_input_payload_stateElements_6;
              buffer_stateElements_7 <= io_input_payload_stateElements_7;
              buffer_stateElements_8 <= io_input_payload_stateElements_8;
              buffer_stateElements_9 <= io_input_payload_stateElements_9;
              buffer_stateElements_10 <= io_input_payload_stateElements_10;
              buffer_stateElements_11 <= io_input_payload_stateElements_11;
            end
          end
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l222) begin
        fsm_counter <= 4'b0000;
      end
    end
  end


endmodule

module StreamArbiter (
  input               io_inputs_0_valid,
  output              io_inputs_0_ready,
  input               io_inputs_0_payload_isFull,
  input      [2:0]    io_inputs_0_payload_fullRound,
  input      [5:0]    io_inputs_0_payload_partialRound,
  input      [3:0]    io_inputs_0_payload_stateSize,
  input      [7:0]    io_inputs_0_payload_stateID,
  input      [254:0]  io_inputs_0_payload_stateElements_0,
  input      [254:0]  io_inputs_0_payload_stateElements_1,
  input      [254:0]  io_inputs_0_payload_stateElements_2,
  input      [254:0]  io_inputs_0_payload_stateElements_3,
  input      [254:0]  io_inputs_0_payload_stateElements_4,
  input      [254:0]  io_inputs_0_payload_stateElements_5,
  input      [254:0]  io_inputs_0_payload_stateElements_6,
  input      [254:0]  io_inputs_0_payload_stateElements_7,
  input      [254:0]  io_inputs_0_payload_stateElements_8,
  input      [254:0]  io_inputs_0_payload_stateElements_9,
  input      [254:0]  io_inputs_0_payload_stateElements_10,
  input      [254:0]  io_inputs_0_payload_stateElements_11,
  input               io_inputs_1_valid,
  output              io_inputs_1_ready,
  input               io_inputs_1_payload_isFull,
  input      [2:0]    io_inputs_1_payload_fullRound,
  input      [5:0]    io_inputs_1_payload_partialRound,
  input      [3:0]    io_inputs_1_payload_stateSize,
  input      [7:0]    io_inputs_1_payload_stateID,
  input      [254:0]  io_inputs_1_payload_stateElements_0,
  input      [254:0]  io_inputs_1_payload_stateElements_1,
  input      [254:0]  io_inputs_1_payload_stateElements_2,
  input      [254:0]  io_inputs_1_payload_stateElements_3,
  input      [254:0]  io_inputs_1_payload_stateElements_4,
  input      [254:0]  io_inputs_1_payload_stateElements_5,
  input      [254:0]  io_inputs_1_payload_stateElements_6,
  input      [254:0]  io_inputs_1_payload_stateElements_7,
  input      [254:0]  io_inputs_1_payload_stateElements_8,
  input      [254:0]  io_inputs_1_payload_stateElements_9,
  input      [254:0]  io_inputs_1_payload_stateElements_10,
  input      [254:0]  io_inputs_1_payload_stateElements_11,
  output              io_output_valid,
  input               io_output_ready,
  output              io_output_payload_isFull,
  output     [2:0]    io_output_payload_fullRound,
  output     [5:0]    io_output_payload_partialRound,
  output     [3:0]    io_output_payload_stateSize,
  output     [7:0]    io_output_payload_stateID,
  output     [254:0]  io_output_payload_stateElements_0,
  output     [254:0]  io_output_payload_stateElements_1,
  output     [254:0]  io_output_payload_stateElements_2,
  output     [254:0]  io_output_payload_stateElements_3,
  output     [254:0]  io_output_payload_stateElements_4,
  output     [254:0]  io_output_payload_stateElements_5,
  output     [254:0]  io_output_payload_stateElements_6,
  output     [254:0]  io_output_payload_stateElements_7,
  output     [254:0]  io_output_payload_stateElements_8,
  output     [254:0]  io_output_payload_stateElements_9,
  output     [254:0]  io_output_payload_stateElements_10,
  output     [254:0]  io_output_payload_stateElements_11,
  output     [0:0]    io_chosen,
  output     [1:0]    io_chosenOH,
  input               clk,
  input               resetn
);

  wire       [1:0]    _zz_maskProposal_1_1;
  wire       [1:0]    _zz_maskProposal_1_2;
  reg                 locked;
  wire                maskProposal_0;
  wire                maskProposal_1;
  reg                 maskLocked_0;
  reg                 maskLocked_1;
  wire                maskRouted_0;
  wire                maskRouted_1;
  wire       [1:0]    _zz_maskProposal_1;
  wire                io_output_fire;
  wire                _zz_io_chosen;

  assign _zz_maskProposal_1_1 = (_zz_maskProposal_1 & (~ _zz_maskProposal_1_2));
  assign _zz_maskProposal_1_2 = (_zz_maskProposal_1 - 2'b01);
  assign maskRouted_0 = (locked ? maskLocked_0 : maskProposal_0);
  assign maskRouted_1 = (locked ? maskLocked_1 : maskProposal_1);
  assign _zz_maskProposal_1 = {io_inputs_1_valid,io_inputs_0_valid};
  assign maskProposal_0 = io_inputs_0_valid;
  assign maskProposal_1 = _zz_maskProposal_1_1[1];
  assign io_output_fire = (io_output_valid && io_output_ready);
  assign io_output_valid = ((io_inputs_0_valid && maskRouted_0) || (io_inputs_1_valid && maskRouted_1));
  assign io_output_payload_isFull = (maskRouted_0 ? io_inputs_0_payload_isFull : io_inputs_1_payload_isFull);
  assign io_output_payload_fullRound = (maskRouted_0 ? io_inputs_0_payload_fullRound : io_inputs_1_payload_fullRound);
  assign io_output_payload_partialRound = (maskRouted_0 ? io_inputs_0_payload_partialRound : io_inputs_1_payload_partialRound);
  assign io_output_payload_stateSize = (maskRouted_0 ? io_inputs_0_payload_stateSize : io_inputs_1_payload_stateSize);
  assign io_output_payload_stateID = (maskRouted_0 ? io_inputs_0_payload_stateID : io_inputs_1_payload_stateID);
  assign io_output_payload_stateElements_0 = (maskRouted_0 ? io_inputs_0_payload_stateElements_0 : io_inputs_1_payload_stateElements_0);
  assign io_output_payload_stateElements_1 = (maskRouted_0 ? io_inputs_0_payload_stateElements_1 : io_inputs_1_payload_stateElements_1);
  assign io_output_payload_stateElements_2 = (maskRouted_0 ? io_inputs_0_payload_stateElements_2 : io_inputs_1_payload_stateElements_2);
  assign io_output_payload_stateElements_3 = (maskRouted_0 ? io_inputs_0_payload_stateElements_3 : io_inputs_1_payload_stateElements_3);
  assign io_output_payload_stateElements_4 = (maskRouted_0 ? io_inputs_0_payload_stateElements_4 : io_inputs_1_payload_stateElements_4);
  assign io_output_payload_stateElements_5 = (maskRouted_0 ? io_inputs_0_payload_stateElements_5 : io_inputs_1_payload_stateElements_5);
  assign io_output_payload_stateElements_6 = (maskRouted_0 ? io_inputs_0_payload_stateElements_6 : io_inputs_1_payload_stateElements_6);
  assign io_output_payload_stateElements_7 = (maskRouted_0 ? io_inputs_0_payload_stateElements_7 : io_inputs_1_payload_stateElements_7);
  assign io_output_payload_stateElements_8 = (maskRouted_0 ? io_inputs_0_payload_stateElements_8 : io_inputs_1_payload_stateElements_8);
  assign io_output_payload_stateElements_9 = (maskRouted_0 ? io_inputs_0_payload_stateElements_9 : io_inputs_1_payload_stateElements_9);
  assign io_output_payload_stateElements_10 = (maskRouted_0 ? io_inputs_0_payload_stateElements_10 : io_inputs_1_payload_stateElements_10);
  assign io_output_payload_stateElements_11 = (maskRouted_0 ? io_inputs_0_payload_stateElements_11 : io_inputs_1_payload_stateElements_11);
  assign io_inputs_0_ready = (maskRouted_0 && io_output_ready);
  assign io_inputs_1_ready = (maskRouted_1 && io_output_ready);
  assign io_chosenOH = {maskRouted_1,maskRouted_0};
  assign _zz_io_chosen = io_chosenOH[1];
  assign io_chosen = _zz_io_chosen;
  always @(posedge clk) begin
    if(!resetn) begin
      locked <= 1'b0;
    end else begin
      if(io_output_valid) begin
        locked <= 1'b1;
      end
      if(io_output_fire) begin
        locked <= 1'b0;
      end
    end
  end

  always @(posedge clk) begin
    if(io_output_valid) begin
      maskLocked_0 <= maskRouted_0;
      maskLocked_1 <= maskRouted_1;
    end
  end


endmodule

module StreamFifo (
  input               io_push_valid,
  output              io_push_ready,
  input               io_push_payload_isFull,
  input      [2:0]    io_push_payload_fullRound,
  input      [5:0]    io_push_payload_partialRound,
  input      [3:0]    io_push_payload_stateSize,
  input      [7:0]    io_push_payload_stateID,
  input      [254:0]  io_push_payload_stateElements_0,
  input      [254:0]  io_push_payload_stateElements_1,
  input      [254:0]  io_push_payload_stateElements_2,
  input      [254:0]  io_push_payload_stateElements_3,
  input      [254:0]  io_push_payload_stateElements_4,
  input      [254:0]  io_push_payload_stateElements_5,
  input      [254:0]  io_push_payload_stateElements_6,
  input      [254:0]  io_push_payload_stateElements_7,
  input      [254:0]  io_push_payload_stateElements_8,
  input      [254:0]  io_push_payload_stateElements_9,
  input      [254:0]  io_push_payload_stateElements_10,
  input      [254:0]  io_push_payload_stateElements_11,
  output              io_pop_valid,
  input               io_pop_ready,
  output              io_pop_payload_isFull,
  output     [2:0]    io_pop_payload_fullRound,
  output     [5:0]    io_pop_payload_partialRound,
  output     [3:0]    io_pop_payload_stateSize,
  output     [7:0]    io_pop_payload_stateID,
  output     [254:0]  io_pop_payload_stateElements_0,
  output     [254:0]  io_pop_payload_stateElements_1,
  output     [254:0]  io_pop_payload_stateElements_2,
  output     [254:0]  io_pop_payload_stateElements_3,
  output     [254:0]  io_pop_payload_stateElements_4,
  output     [254:0]  io_pop_payload_stateElements_5,
  output     [254:0]  io_pop_payload_stateElements_6,
  output     [254:0]  io_pop_payload_stateElements_7,
  output     [254:0]  io_pop_payload_stateElements_8,
  output     [254:0]  io_pop_payload_stateElements_9,
  output     [254:0]  io_pop_payload_stateElements_10,
  output     [254:0]  io_pop_payload_stateElements_11,
  input               io_flush,
  output     [8:0]    io_occupancy,
  output     [8:0]    io_availability,
  input               clk,
  input               resetn
);

  reg        [3081:0] _zz_logic_ram_port0;
  wire       [7:0]    _zz_logic_pushPtr_valueNext;
  wire       [0:0]    _zz_logic_pushPtr_valueNext_1;
  wire       [7:0]    _zz_logic_popPtr_valueNext;
  wire       [0:0]    _zz_logic_popPtr_valueNext_1;
  wire                _zz_logic_ram_port;
  wire                _zz__zz_io_pop_payload_isFull;
  wire       [3081:0] _zz_logic_ram_port_1;
  wire       [7:0]    _zz_io_availability;
  reg                 _zz_1;
  reg                 logic_pushPtr_willIncrement;
  reg                 logic_pushPtr_willClear;
  reg        [7:0]    logic_pushPtr_valueNext;
  reg        [7:0]    logic_pushPtr_value;
  wire                logic_pushPtr_willOverflowIfInc;
  wire                logic_pushPtr_willOverflow;
  reg                 logic_popPtr_willIncrement;
  reg                 logic_popPtr_willClear;
  reg        [7:0]    logic_popPtr_valueNext;
  reg        [7:0]    logic_popPtr_value;
  wire                logic_popPtr_willOverflowIfInc;
  wire                logic_popPtr_willOverflow;
  wire                logic_ptrMatch;
  reg                 logic_risingOccupancy;
  wire                logic_pushing;
  wire                logic_popping;
  wire                logic_empty;
  wire                logic_full;
  reg                 _zz_io_pop_valid;
  wire       [3081:0] _zz_io_pop_payload_isFull;
  wire       [3059:0] _zz_io_pop_payload_stateElements_0;
  wire                when_Stream_l954;
  wire       [7:0]    logic_ptrDif;
  reg [3081:0] logic_ram [0:255];

  assign _zz_logic_pushPtr_valueNext_1 = logic_pushPtr_willIncrement;
  assign _zz_logic_pushPtr_valueNext = {7'd0, _zz_logic_pushPtr_valueNext_1};
  assign _zz_logic_popPtr_valueNext_1 = logic_popPtr_willIncrement;
  assign _zz_logic_popPtr_valueNext = {7'd0, _zz_logic_popPtr_valueNext_1};
  assign _zz_io_availability = (logic_popPtr_value - logic_pushPtr_value);
  assign _zz__zz_io_pop_payload_isFull = 1'b1;
  assign _zz_logic_ram_port_1 = {{io_push_payload_stateElements_11,{io_push_payload_stateElements_10,{io_push_payload_stateElements_9,{io_push_payload_stateElements_8,{io_push_payload_stateElements_7,{io_push_payload_stateElements_6,{io_push_payload_stateElements_5,{io_push_payload_stateElements_4,{io_push_payload_stateElements_3,{io_push_payload_stateElements_2,{io_push_payload_stateElements_1,io_push_payload_stateElements_0}}}}}}}}}}},{io_push_payload_stateID,{io_push_payload_stateSize,{io_push_payload_partialRound,{io_push_payload_fullRound,io_push_payload_isFull}}}}};
  always @(posedge clk) begin
    if(_zz__zz_io_pop_payload_isFull) begin
      _zz_logic_ram_port0 <= logic_ram[logic_popPtr_valueNext];
    end
  end

  always @(posedge clk) begin
    if(_zz_1) begin
      logic_ram[logic_pushPtr_value] <= _zz_logic_ram_port_1;
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(logic_pushing) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willIncrement = 1'b0;
    if(logic_pushing) begin
      logic_pushPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_pushPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_pushPtr_willClear = 1'b1;
    end
  end

  assign logic_pushPtr_willOverflowIfInc = (logic_pushPtr_value == 8'hff);
  assign logic_pushPtr_willOverflow = (logic_pushPtr_willOverflowIfInc && logic_pushPtr_willIncrement);
  always @(*) begin
    logic_pushPtr_valueNext = (logic_pushPtr_value + _zz_logic_pushPtr_valueNext);
    if(logic_pushPtr_willClear) begin
      logic_pushPtr_valueNext = 8'h0;
    end
  end

  always @(*) begin
    logic_popPtr_willIncrement = 1'b0;
    if(logic_popping) begin
      logic_popPtr_willIncrement = 1'b1;
    end
  end

  always @(*) begin
    logic_popPtr_willClear = 1'b0;
    if(io_flush) begin
      logic_popPtr_willClear = 1'b1;
    end
  end

  assign logic_popPtr_willOverflowIfInc = (logic_popPtr_value == 8'hff);
  assign logic_popPtr_willOverflow = (logic_popPtr_willOverflowIfInc && logic_popPtr_willIncrement);
  always @(*) begin
    logic_popPtr_valueNext = (logic_popPtr_value + _zz_logic_popPtr_valueNext);
    if(logic_popPtr_willClear) begin
      logic_popPtr_valueNext = 8'h0;
    end
  end

  assign logic_ptrMatch = (logic_pushPtr_value == logic_popPtr_value);
  assign logic_pushing = (io_push_valid && io_push_ready);
  assign logic_popping = (io_pop_valid && io_pop_ready);
  assign logic_empty = (logic_ptrMatch && (! logic_risingOccupancy));
  assign logic_full = (logic_ptrMatch && logic_risingOccupancy);
  assign io_push_ready = (! logic_full);
  assign io_pop_valid = ((! logic_empty) && (! (_zz_io_pop_valid && (! logic_full))));
  assign _zz_io_pop_payload_isFull = _zz_logic_ram_port0;
  assign _zz_io_pop_payload_stateElements_0 = _zz_io_pop_payload_isFull[3081 : 22];
  assign io_pop_payload_isFull = _zz_io_pop_payload_isFull[0];
  assign io_pop_payload_fullRound = _zz_io_pop_payload_isFull[3 : 1];
  assign io_pop_payload_partialRound = _zz_io_pop_payload_isFull[9 : 4];
  assign io_pop_payload_stateSize = _zz_io_pop_payload_isFull[13 : 10];
  assign io_pop_payload_stateID = _zz_io_pop_payload_isFull[21 : 14];
  assign io_pop_payload_stateElements_0 = _zz_io_pop_payload_stateElements_0[254 : 0];
  assign io_pop_payload_stateElements_1 = _zz_io_pop_payload_stateElements_0[509 : 255];
  assign io_pop_payload_stateElements_2 = _zz_io_pop_payload_stateElements_0[764 : 510];
  assign io_pop_payload_stateElements_3 = _zz_io_pop_payload_stateElements_0[1019 : 765];
  assign io_pop_payload_stateElements_4 = _zz_io_pop_payload_stateElements_0[1274 : 1020];
  assign io_pop_payload_stateElements_5 = _zz_io_pop_payload_stateElements_0[1529 : 1275];
  assign io_pop_payload_stateElements_6 = _zz_io_pop_payload_stateElements_0[1784 : 1530];
  assign io_pop_payload_stateElements_7 = _zz_io_pop_payload_stateElements_0[2039 : 1785];
  assign io_pop_payload_stateElements_8 = _zz_io_pop_payload_stateElements_0[2294 : 2040];
  assign io_pop_payload_stateElements_9 = _zz_io_pop_payload_stateElements_0[2549 : 2295];
  assign io_pop_payload_stateElements_10 = _zz_io_pop_payload_stateElements_0[2804 : 2550];
  assign io_pop_payload_stateElements_11 = _zz_io_pop_payload_stateElements_0[3059 : 2805];
  assign when_Stream_l954 = (logic_pushing != logic_popping);
  assign logic_ptrDif = (logic_pushPtr_value - logic_popPtr_value);
  assign io_occupancy = {(logic_risingOccupancy && logic_ptrMatch),logic_ptrDif};
  assign io_availability = {((! logic_risingOccupancy) && logic_ptrMatch),_zz_io_availability};
  always @(posedge clk) begin
    if(!resetn) begin
      logic_pushPtr_value <= 8'h0;
      logic_popPtr_value <= 8'h0;
      logic_risingOccupancy <= 1'b0;
      _zz_io_pop_valid <= 1'b0;
    end else begin
      logic_pushPtr_value <= logic_pushPtr_valueNext;
      logic_popPtr_value <= logic_popPtr_valueNext;
      _zz_io_pop_valid <= (logic_popPtr_valueNext == logic_pushPtr_value);
      if(when_Stream_l954) begin
        logic_risingOccupancy <= logic_pushing;
      end
      if(io_flush) begin
        logic_risingOccupancy <= 1'b0;
      end
    end
  end


endmodule

module StreamDemux (
  input      [0:0]    io_select,
  input               io_input_valid,
  output reg          io_input_ready,
  input               io_input_payload_isFull,
  input      [2:0]    io_input_payload_fullRound,
  input      [5:0]    io_input_payload_partialRound,
  input      [3:0]    io_input_payload_stateSize,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElements_0,
  input      [254:0]  io_input_payload_stateElements_1,
  input      [254:0]  io_input_payload_stateElements_2,
  input      [254:0]  io_input_payload_stateElements_3,
  input      [254:0]  io_input_payload_stateElements_4,
  input      [254:0]  io_input_payload_stateElements_5,
  input      [254:0]  io_input_payload_stateElements_6,
  input      [254:0]  io_input_payload_stateElements_7,
  input      [254:0]  io_input_payload_stateElements_8,
  input      [254:0]  io_input_payload_stateElements_9,
  input      [254:0]  io_input_payload_stateElements_10,
  input      [254:0]  io_input_payload_stateElements_11,
  output reg          io_outputs_0_valid,
  input               io_outputs_0_ready,
  output              io_outputs_0_payload_isFull,
  output     [2:0]    io_outputs_0_payload_fullRound,
  output     [5:0]    io_outputs_0_payload_partialRound,
  output     [3:0]    io_outputs_0_payload_stateSize,
  output     [7:0]    io_outputs_0_payload_stateID,
  output     [254:0]  io_outputs_0_payload_stateElements_0,
  output     [254:0]  io_outputs_0_payload_stateElements_1,
  output     [254:0]  io_outputs_0_payload_stateElements_2,
  output     [254:0]  io_outputs_0_payload_stateElements_3,
  output     [254:0]  io_outputs_0_payload_stateElements_4,
  output     [254:0]  io_outputs_0_payload_stateElements_5,
  output     [254:0]  io_outputs_0_payload_stateElements_6,
  output     [254:0]  io_outputs_0_payload_stateElements_7,
  output     [254:0]  io_outputs_0_payload_stateElements_8,
  output     [254:0]  io_outputs_0_payload_stateElements_9,
  output     [254:0]  io_outputs_0_payload_stateElements_10,
  output     [254:0]  io_outputs_0_payload_stateElements_11,
  output reg          io_outputs_1_valid,
  input               io_outputs_1_ready,
  output              io_outputs_1_payload_isFull,
  output     [2:0]    io_outputs_1_payload_fullRound,
  output     [5:0]    io_outputs_1_payload_partialRound,
  output     [3:0]    io_outputs_1_payload_stateSize,
  output     [7:0]    io_outputs_1_payload_stateID,
  output     [254:0]  io_outputs_1_payload_stateElements_0,
  output     [254:0]  io_outputs_1_payload_stateElements_1,
  output     [254:0]  io_outputs_1_payload_stateElements_2,
  output     [254:0]  io_outputs_1_payload_stateElements_3,
  output     [254:0]  io_outputs_1_payload_stateElements_4,
  output     [254:0]  io_outputs_1_payload_stateElements_5,
  output     [254:0]  io_outputs_1_payload_stateElements_6,
  output     [254:0]  io_outputs_1_payload_stateElements_7,
  output     [254:0]  io_outputs_1_payload_stateElements_8,
  output     [254:0]  io_outputs_1_payload_stateElements_9,
  output     [254:0]  io_outputs_1_payload_stateElements_10,
  output     [254:0]  io_outputs_1_payload_stateElements_11
);

  wire                when_Stream_l764;
  wire                when_Stream_l764_1;

  always @(*) begin
    io_input_ready = 1'b0;
    if(!when_Stream_l764) begin
      io_input_ready = io_outputs_0_ready;
    end
    if(!when_Stream_l764_1) begin
      io_input_ready = io_outputs_1_ready;
    end
  end

  assign io_outputs_0_payload_isFull = io_input_payload_isFull;
  assign io_outputs_0_payload_fullRound = io_input_payload_fullRound;
  assign io_outputs_0_payload_partialRound = io_input_payload_partialRound;
  assign io_outputs_0_payload_stateSize = io_input_payload_stateSize;
  assign io_outputs_0_payload_stateID = io_input_payload_stateID;
  assign io_outputs_0_payload_stateElements_0 = io_input_payload_stateElements_0;
  assign io_outputs_0_payload_stateElements_1 = io_input_payload_stateElements_1;
  assign io_outputs_0_payload_stateElements_2 = io_input_payload_stateElements_2;
  assign io_outputs_0_payload_stateElements_3 = io_input_payload_stateElements_3;
  assign io_outputs_0_payload_stateElements_4 = io_input_payload_stateElements_4;
  assign io_outputs_0_payload_stateElements_5 = io_input_payload_stateElements_5;
  assign io_outputs_0_payload_stateElements_6 = io_input_payload_stateElements_6;
  assign io_outputs_0_payload_stateElements_7 = io_input_payload_stateElements_7;
  assign io_outputs_0_payload_stateElements_8 = io_input_payload_stateElements_8;
  assign io_outputs_0_payload_stateElements_9 = io_input_payload_stateElements_9;
  assign io_outputs_0_payload_stateElements_10 = io_input_payload_stateElements_10;
  assign io_outputs_0_payload_stateElements_11 = io_input_payload_stateElements_11;
  assign when_Stream_l764 = (1'b0 != io_select);
  always @(*) begin
    if(when_Stream_l764) begin
      io_outputs_0_valid = 1'b0;
    end else begin
      io_outputs_0_valid = io_input_valid;
    end
  end

  assign io_outputs_1_payload_isFull = io_input_payload_isFull;
  assign io_outputs_1_payload_fullRound = io_input_payload_fullRound;
  assign io_outputs_1_payload_partialRound = io_input_payload_partialRound;
  assign io_outputs_1_payload_stateSize = io_input_payload_stateSize;
  assign io_outputs_1_payload_stateID = io_input_payload_stateID;
  assign io_outputs_1_payload_stateElements_0 = io_input_payload_stateElements_0;
  assign io_outputs_1_payload_stateElements_1 = io_input_payload_stateElements_1;
  assign io_outputs_1_payload_stateElements_2 = io_input_payload_stateElements_2;
  assign io_outputs_1_payload_stateElements_3 = io_input_payload_stateElements_3;
  assign io_outputs_1_payload_stateElements_4 = io_input_payload_stateElements_4;
  assign io_outputs_1_payload_stateElements_5 = io_input_payload_stateElements_5;
  assign io_outputs_1_payload_stateElements_6 = io_input_payload_stateElements_6;
  assign io_outputs_1_payload_stateElements_7 = io_input_payload_stateElements_7;
  assign io_outputs_1_payload_stateElements_8 = io_input_payload_stateElements_8;
  assign io_outputs_1_payload_stateElements_9 = io_input_payload_stateElements_9;
  assign io_outputs_1_payload_stateElements_10 = io_input_payload_stateElements_10;
  assign io_outputs_1_payload_stateElements_11 = io_input_payload_stateElements_11;
  assign when_Stream_l764_1 = (1'b1 != io_select);
  always @(*) begin
    if(when_Stream_l764_1) begin
      io_outputs_1_valid = 1'b0;
    end else begin
      io_outputs_1_valid = io_input_valid;
    end
  end


endmodule

module MDSMatrixAdders (
  input               io_input_valid,
  input               io_input_payload_isFull,
  input      [2:0]    io_input_payload_fullRound,
  input      [5:0]    io_input_payload_partialRound,
  input      [3:0]    io_input_payload_stateSize,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElements_0,
  input      [254:0]  io_input_payload_stateElements_1,
  input      [254:0]  io_input_payload_stateElements_2,
  input      [254:0]  io_input_payload_stateElements_3,
  input      [254:0]  io_input_payload_stateElements_4,
  input      [254:0]  io_input_payload_stateElements_5,
  input      [254:0]  io_input_payload_stateElements_6,
  input      [254:0]  io_input_payload_stateElements_7,
  input      [254:0]  io_input_payload_stateElements_8,
  input      [254:0]  io_input_payload_stateElements_9,
  input      [254:0]  io_input_payload_stateElements_10,
  input      [254:0]  io_input_payload_stateElements_11,
  output reg          io_output_valid,
  output reg          io_output_payload_isFull,
  output reg [2:0]    io_output_payload_fullRound,
  output reg [5:0]    io_output_payload_partialRound,
  output reg [3:0]    io_output_payload_stateSize,
  output reg [7:0]    io_output_payload_stateID,
  output reg [254:0]  io_output_payload_stateElements_0,
  output reg [254:0]  io_output_payload_stateElements_1,
  output reg [254:0]  io_output_payload_stateElements_2,
  output reg [254:0]  io_output_payload_stateElements_3,
  output reg [254:0]  io_output_payload_stateElements_4,
  output reg [254:0]  io_output_payload_stateElements_5,
  output reg [254:0]  io_output_payload_stateElements_6,
  output reg [254:0]  io_output_payload_stateElements_7,
  output reg [254:0]  io_output_payload_stateElements_8,
  output reg [254:0]  io_output_payload_stateElements_9,
  output reg [254:0]  io_output_payload_stateElements_10,
  output reg [254:0]  io_output_payload_stateElements_11,
  input               clk,
  input               resetn
);
  localparam fullRound_deserialization_enumDef_BOOT = 2'd0;
  localparam fullRound_deserialization_enumDef_IDLE = 2'd1;
  localparam fullRound_deserialization_enumDef_BUSY = 2'd2;
  localparam fullRound_deserialization_enumDef_DONE = 2'd3;

  reg                 adderTree_1_io_input_valid;
  reg        [254:0]  adderTree_1_io_input_payload_0;
  reg        [254:0]  adderTree_1_io_input_payload_1;
  reg        [254:0]  adderTree_1_io_input_payload_2;
  reg        [254:0]  adderTree_1_io_input_payload_3;
  reg        [254:0]  adderTree_1_io_input_payload_4;
  reg        [254:0]  adderTree_1_io_input_payload_5;
  reg        [254:0]  adderTree_1_io_input_payload_6;
  reg        [254:0]  adderTree_1_io_input_payload_7;
  reg        [254:0]  adderTree_1_io_input_payload_8;
  reg        [254:0]  adderTree_1_io_input_payload_9;
  reg        [254:0]  adderTree_1_io_input_payload_10;
  reg        [254:0]  adderTree_1_io_input_payload_11;
  wire                adderTree_1_io_output_valid;
  wire       [254:0]  adderTree_1_io_output_payload;
  wire                fullRound_shiftMat_io_output_valid;
  wire                fullRound_shiftMat_io_output_payload_isFull;
  wire       [2:0]    fullRound_shiftMat_io_output_payload_fullRound;
  wire       [5:0]    fullRound_shiftMat_io_output_payload_partialRound;
  wire       [3:0]    fullRound_shiftMat_io_output_payload_stateSize;
  wire       [7:0]    fullRound_shiftMat_io_output_payload_stateID;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_0;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_1;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_2;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_3;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_4;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_5;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_6;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_7;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_8;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_9;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_10;
  wire       [254:0]  fullRound_shiftMat_io_output_payload_stateElements_11;
  reg                 _zz_partialRound_bufferOutMuxed_valid_3;
  reg                 _zz_partialRound_bufferOutMuxed_payload_isFull;
  reg        [2:0]    _zz_partialRound_bufferOutMuxed_payload_fullRound;
  reg        [5:0]    _zz_partialRound_bufferOutMuxed_payload_partialRound;
  reg        [3:0]    _zz_partialRound_bufferOutMuxed_payload_stateSize;
  reg        [7:0]    _zz_partialRound_bufferOutMuxed_payload_stateID;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_0;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_1;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_2;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_3;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_4;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_5;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_6;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_7;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_8;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_9;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_10;
  reg        [254:0]  _zz_partialRound_bufferOutMuxed_payload_stateElements_11;
  wire       [3:0]    _zz_when_MDSMatrixAdders_l147;
  wire                partialRound_input_valid;
  wire                partialRound_input_payload_isFull;
  wire       [2:0]    partialRound_input_payload_fullRound;
  wire       [5:0]    partialRound_input_payload_partialRound;
  wire       [3:0]    partialRound_input_payload_stateSize;
  wire       [7:0]    partialRound_input_payload_stateID;
  wire       [254:0]  partialRound_input_payload_stateElements_0;
  wire       [254:0]  partialRound_input_payload_stateElements_1;
  wire       [254:0]  partialRound_input_payload_stateElements_2;
  wire       [254:0]  partialRound_input_payload_stateElements_3;
  wire       [254:0]  partialRound_input_payload_stateElements_4;
  wire       [254:0]  partialRound_input_payload_stateElements_5;
  wire       [254:0]  partialRound_input_payload_stateElements_6;
  wire       [254:0]  partialRound_input_payload_stateElements_7;
  wire       [254:0]  partialRound_input_payload_stateElements_8;
  wire       [254:0]  partialRound_input_payload_stateElements_9;
  wire       [254:0]  partialRound_input_payload_stateElements_10;
  wire       [254:0]  partialRound_input_payload_stateElements_11;
  wire                partialRound_inputBuffered_0_valid;
  wire                partialRound_inputBuffered_0_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_0_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_0_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_0_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_0_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_0_payload_stateElements_11;
  wire                partialRound_inputBuffered_1_valid;
  wire                partialRound_inputBuffered_1_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_1_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_1_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_1_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_1_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_1_payload_stateElements_11;
  wire                partialRound_inputBuffered_2_valid;
  wire                partialRound_inputBuffered_2_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_2_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_2_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_2_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_2_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_2_payload_stateElements_11;
  wire                partialRound_inputBuffered_3_valid;
  wire                partialRound_inputBuffered_3_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_3_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_3_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_3_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_3_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_3_payload_stateElements_11;
  wire                partialRound_inputBuffered_4_valid;
  wire                partialRound_inputBuffered_4_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_4_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_4_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_4_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_4_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_4_payload_stateElements_11;
  wire                partialRound_inputBuffered_5_valid;
  wire                partialRound_inputBuffered_5_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_5_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_5_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_5_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_5_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_5_payload_stateElements_11;
  wire                partialRound_inputBuffered_6_valid;
  wire                partialRound_inputBuffered_6_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_6_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_6_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_6_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_6_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_6_payload_stateElements_11;
  wire                partialRound_inputBuffered_7_valid;
  wire                partialRound_inputBuffered_7_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_7_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_7_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_7_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_7_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_7_payload_stateElements_11;
  wire                partialRound_inputBuffered_8_valid;
  wire                partialRound_inputBuffered_8_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_8_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_8_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_8_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_8_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_8_payload_stateElements_11;
  wire                partialRound_inputBuffered_9_valid;
  wire                partialRound_inputBuffered_9_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_9_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_9_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_9_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_9_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_9_payload_stateElements_11;
  wire                partialRound_inputBuffered_10_valid;
  wire                partialRound_inputBuffered_10_payload_isFull;
  wire       [2:0]    partialRound_inputBuffered_10_payload_fullRound;
  wire       [5:0]    partialRound_inputBuffered_10_payload_partialRound;
  wire       [3:0]    partialRound_inputBuffered_10_payload_stateSize;
  wire       [7:0]    partialRound_inputBuffered_10_payload_stateID;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_0;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_1;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_2;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_3;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_4;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_5;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_6;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_7;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_8;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_9;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_10;
  wire       [254:0]  partialRound_inputBuffered_10_payload_stateElements_11;
  reg                 partialRound_input_regNext_valid;
  reg                 partialRound_input_regNext_payload_isFull;
  reg        [2:0]    partialRound_input_regNext_payload_fullRound;
  reg        [5:0]    partialRound_input_regNext_payload_partialRound;
  reg        [3:0]    partialRound_input_regNext_payload_stateSize;
  reg        [7:0]    partialRound_input_regNext_payload_stateID;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_input_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_0_regNext_valid;
  reg                 partialRound_inputBuffered_0_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_0_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_0_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_0_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_0_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_0_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_1_regNext_valid;
  reg                 partialRound_inputBuffered_1_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_1_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_1_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_1_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_1_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_1_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_2_regNext_valid;
  reg                 partialRound_inputBuffered_2_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_2_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_2_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_2_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_2_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_2_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_3_regNext_valid;
  reg                 partialRound_inputBuffered_3_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_3_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_3_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_3_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_3_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_3_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_4_regNext_valid;
  reg                 partialRound_inputBuffered_4_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_4_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_4_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_4_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_4_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_4_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_5_regNext_valid;
  reg                 partialRound_inputBuffered_5_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_5_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_5_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_5_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_5_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_5_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_6_regNext_valid;
  reg                 partialRound_inputBuffered_6_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_6_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_6_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_6_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_6_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_6_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_7_regNext_valid;
  reg                 partialRound_inputBuffered_7_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_7_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_7_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_7_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_7_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_7_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_8_regNext_valid;
  reg                 partialRound_inputBuffered_8_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_8_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_8_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_8_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_8_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_8_regNext_payload_stateElements_11;
  reg                 partialRound_inputBuffered_9_regNext_valid;
  reg                 partialRound_inputBuffered_9_regNext_payload_isFull;
  reg        [2:0]    partialRound_inputBuffered_9_regNext_payload_fullRound;
  reg        [5:0]    partialRound_inputBuffered_9_regNext_payload_partialRound;
  reg        [3:0]    partialRound_inputBuffered_9_regNext_payload_stateSize;
  reg        [7:0]    partialRound_inputBuffered_9_regNext_payload_stateID;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_0;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_1;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_2;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_3;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_4;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_5;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_6;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_7;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_8;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_9;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_10;
  reg        [254:0]  partialRound_inputBuffered_9_regNext_payload_stateElements_11;
  wire                partialRound_bufferOut_0_valid;
  wire                partialRound_bufferOut_0_payload_isFull;
  wire       [2:0]    partialRound_bufferOut_0_payload_fullRound;
  wire       [5:0]    partialRound_bufferOut_0_payload_partialRound;
  wire       [3:0]    partialRound_bufferOut_0_payload_stateSize;
  wire       [7:0]    partialRound_bufferOut_0_payload_stateID;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_0;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_1;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_2;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_3;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_4;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_5;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_6;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_7;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_8;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_9;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_10;
  wire       [254:0]  partialRound_bufferOut_0_payload_stateElements_11;
  wire                partialRound_bufferOut_1_valid;
  wire                partialRound_bufferOut_1_payload_isFull;
  wire       [2:0]    partialRound_bufferOut_1_payload_fullRound;
  wire       [5:0]    partialRound_bufferOut_1_payload_partialRound;
  wire       [3:0]    partialRound_bufferOut_1_payload_stateSize;
  wire       [7:0]    partialRound_bufferOut_1_payload_stateID;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_0;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_1;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_2;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_3;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_4;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_5;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_6;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_7;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_8;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_9;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_10;
  wire       [254:0]  partialRound_bufferOut_1_payload_stateElements_11;
  wire                partialRound_bufferOut_2_valid;
  wire                partialRound_bufferOut_2_payload_isFull;
  wire       [2:0]    partialRound_bufferOut_2_payload_fullRound;
  wire       [5:0]    partialRound_bufferOut_2_payload_partialRound;
  wire       [3:0]    partialRound_bufferOut_2_payload_stateSize;
  wire       [7:0]    partialRound_bufferOut_2_payload_stateID;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_0;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_1;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_2;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_3;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_4;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_5;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_6;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_7;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_8;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_9;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_10;
  wire       [254:0]  partialRound_bufferOut_2_payload_stateElements_11;
  wire                partialRound_bufferOut_3_valid;
  wire                partialRound_bufferOut_3_payload_isFull;
  wire       [2:0]    partialRound_bufferOut_3_payload_fullRound;
  wire       [5:0]    partialRound_bufferOut_3_payload_partialRound;
  wire       [3:0]    partialRound_bufferOut_3_payload_stateSize;
  wire       [7:0]    partialRound_bufferOut_3_payload_stateID;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_0;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_1;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_2;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_3;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_4;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_5;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_6;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_7;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_8;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_9;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_10;
  wire       [254:0]  partialRound_bufferOut_3_payload_stateElements_11;
  wire                _zz_partialRound_bufferOutMuxed_valid;
  wire                _zz_partialRound_bufferOutMuxed_valid_1;
  wire       [1:0]    _zz_partialRound_bufferOutMuxed_valid_2;
  wire                partialRound_bufferOutMuxed_valid;
  wire                partialRound_bufferOutMuxed_payload_isFull;
  wire       [2:0]    partialRound_bufferOutMuxed_payload_fullRound;
  wire       [5:0]    partialRound_bufferOutMuxed_payload_partialRound;
  wire       [3:0]    partialRound_bufferOutMuxed_payload_stateSize;
  wire       [7:0]    partialRound_bufferOutMuxed_payload_stateID;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_0;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_1;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_2;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_3;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_4;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_5;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_6;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_7;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_8;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_9;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_10;
  wire       [254:0]  partialRound_bufferOutMuxed_payload_stateElements_11;
  reg                 partialRound_partialFlag;
  wire                when_MDSMatrixAdders_l67;
  wire                partialRound_bufferOutMuxed_takeWhen_valid;
  wire                partialRound_bufferOutMuxed_takeWhen_payload_isFull;
  wire       [2:0]    partialRound_bufferOutMuxed_takeWhen_payload_fullRound;
  wire       [5:0]    partialRound_bufferOutMuxed_takeWhen_payload_partialRound;
  wire       [3:0]    partialRound_bufferOutMuxed_takeWhen_payload_stateSize;
  wire       [7:0]    partialRound_bufferOutMuxed_takeWhen_payload_stateID;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_0;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_1;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_2;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_3;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_4;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_5;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_6;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_7;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_8;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_9;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_10;
  wire       [254:0]  partialRound_bufferOutMuxed_takeWhen_payload_stateElements_11;
  reg                 partialRound_tempInput_valid;
  reg                 partialRound_tempInput_payload_isFull;
  reg        [2:0]    partialRound_tempInput_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_payload_stateID;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_payload_stateElements_11;
  reg        [254:0]  _zz_partialRound_adderTreeInput_payload_1;
  reg        [254:0]  _zz_partialRound_adderTreeInput_payload_2;
  reg        [254:0]  _zz_partialRound_adderTreeInput_payload_3;
  reg        [254:0]  _zz_partialRound_adderTreeInput_payload_4;
  wire                when_MDSMatrixAdders_l75;
  wire                when_MDSMatrixAdders_l77;
  wire                partialRound_adderTreeInput_valid;
  wire       [254:0]  partialRound_adderTreeInput_payload_0;
  wire       [254:0]  partialRound_adderTreeInput_payload_1;
  wire       [254:0]  partialRound_adderTreeInput_payload_2;
  wire       [254:0]  partialRound_adderTreeInput_payload_3;
  wire       [254:0]  partialRound_adderTreeInput_payload_4;
  wire       [254:0]  partialRound_adderTreeInput_payload_5;
  wire       [254:0]  partialRound_adderTreeInput_payload_6;
  wire       [254:0]  partialRound_adderTreeInput_payload_7;
  wire       [254:0]  partialRound_adderTreeInput_payload_8;
  wire       [254:0]  partialRound_adderTreeInput_payload_9;
  wire       [254:0]  partialRound_adderTreeInput_payload_10;
  wire       [254:0]  partialRound_adderTreeInput_payload_11;
  reg                 partialRound_tempInput_delay_1_valid;
  reg                 partialRound_tempInput_delay_1_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_1_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_1_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_1_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_1_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_1_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_2_valid;
  reg                 partialRound_tempInput_delay_2_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_2_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_2_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_2_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_2_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_2_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_3_valid;
  reg                 partialRound_tempInput_delay_3_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_3_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_3_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_3_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_3_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_3_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_4_valid;
  reg                 partialRound_tempInput_delay_4_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_4_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_4_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_4_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_4_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_4_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_5_valid;
  reg                 partialRound_tempInput_delay_5_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_5_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_5_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_5_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_5_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_5_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_6_valid;
  reg                 partialRound_tempInput_delay_6_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_6_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_6_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_6_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_6_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_6_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_7_valid;
  reg                 partialRound_tempInput_delay_7_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_7_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_7_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_7_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_7_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_7_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_8_valid;
  reg                 partialRound_tempInput_delay_8_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_8_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_8_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_8_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_8_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_8_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_9_valid;
  reg                 partialRound_tempInput_delay_9_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_9_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_9_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_9_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_9_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_9_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_10_valid;
  reg                 partialRound_tempInput_delay_10_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_10_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_10_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_10_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_10_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_10_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_11_valid;
  reg                 partialRound_tempInput_delay_11_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_11_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_11_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_11_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_11_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_11_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_12_valid;
  reg                 partialRound_tempInput_delay_12_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_12_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_12_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_12_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_12_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_12_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_13_valid;
  reg                 partialRound_tempInput_delay_13_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_13_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_13_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_13_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_13_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_13_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_14_valid;
  reg                 partialRound_tempInput_delay_14_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_14_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_14_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_14_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_14_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_14_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_15_valid;
  reg                 partialRound_tempInput_delay_15_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_15_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_15_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_15_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_15_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_15_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_16_valid;
  reg                 partialRound_tempInput_delay_16_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_16_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_16_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_16_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_16_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_16_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_17_valid;
  reg                 partialRound_tempInput_delay_17_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_17_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_17_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_17_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_17_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_17_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_18_valid;
  reg                 partialRound_tempInput_delay_18_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_18_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_18_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_18_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_18_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_18_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_19_valid;
  reg                 partialRound_tempInput_delay_19_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_19_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_19_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_19_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_19_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_19_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_20_valid;
  reg                 partialRound_tempInput_delay_20_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_20_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_20_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_20_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_20_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_20_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_21_valid;
  reg                 partialRound_tempInput_delay_21_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_21_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_21_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_21_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_21_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_21_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_22_valid;
  reg                 partialRound_tempInput_delay_22_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_22_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_22_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_22_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_22_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_22_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_23_valid;
  reg                 partialRound_tempInput_delay_23_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_23_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_23_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_23_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_23_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_23_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_24_valid;
  reg                 partialRound_tempInput_delay_24_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_24_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_24_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_24_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_24_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_24_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_25_valid;
  reg                 partialRound_tempInput_delay_25_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_25_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_25_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_25_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_25_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_25_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_26_valid;
  reg                 partialRound_tempInput_delay_26_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_26_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_26_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_26_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_26_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_26_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_27_valid;
  reg                 partialRound_tempInput_delay_27_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_27_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_27_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_27_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_27_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_27_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_28_valid;
  reg                 partialRound_tempInput_delay_28_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_28_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_28_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_28_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_28_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_28_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_29_valid;
  reg                 partialRound_tempInput_delay_29_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_29_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_29_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_29_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_29_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_29_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_30_valid;
  reg                 partialRound_tempInput_delay_30_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_30_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_30_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_30_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_30_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_30_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_31_valid;
  reg                 partialRound_tempInput_delay_31_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_31_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_31_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_31_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_31_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_31_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_32_valid;
  reg                 partialRound_tempInput_delay_32_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_32_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_32_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_32_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_32_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_32_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_33_valid;
  reg                 partialRound_tempInput_delay_33_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_33_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_33_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_33_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_33_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_33_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_34_valid;
  reg                 partialRound_tempInput_delay_34_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_34_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_34_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_34_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_34_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_34_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_35_valid;
  reg                 partialRound_tempInput_delay_35_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_35_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_35_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_35_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_35_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_35_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_36_valid;
  reg                 partialRound_tempInput_delay_36_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_36_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_36_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_36_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_36_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_36_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_37_valid;
  reg                 partialRound_tempInput_delay_37_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_37_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_37_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_37_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_37_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_37_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_38_valid;
  reg                 partialRound_tempInput_delay_38_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_38_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_38_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_38_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_38_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_38_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_39_valid;
  reg                 partialRound_tempInput_delay_39_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_39_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_39_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_39_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_39_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_39_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_40_valid;
  reg                 partialRound_tempInput_delay_40_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_40_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_40_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_40_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_40_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_40_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_41_valid;
  reg                 partialRound_tempInput_delay_41_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_41_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_41_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_41_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_41_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_41_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_42_valid;
  reg                 partialRound_tempInput_delay_42_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_42_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_42_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_42_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_42_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_42_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_43_valid;
  reg                 partialRound_tempInput_delay_43_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_43_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_43_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_43_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_43_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_43_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_44_valid;
  reg                 partialRound_tempInput_delay_44_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_44_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_44_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_44_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_44_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_44_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_45_valid;
  reg                 partialRound_tempInput_delay_45_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_45_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_45_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_45_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_45_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_45_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_46_valid;
  reg                 partialRound_tempInput_delay_46_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_46_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_46_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_46_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_46_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_46_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_47_valid;
  reg                 partialRound_tempInput_delay_47_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_47_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_47_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_47_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_47_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_47_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_48_valid;
  reg                 partialRound_tempInput_delay_48_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_48_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_48_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_48_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_48_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_48_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_49_valid;
  reg                 partialRound_tempInput_delay_49_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_49_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_49_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_49_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_49_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_49_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_50_valid;
  reg                 partialRound_tempInput_delay_50_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_50_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_50_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_50_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_50_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_50_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_51_valid;
  reg                 partialRound_tempInput_delay_51_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_51_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_51_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_51_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_51_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_51_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_52_valid;
  reg                 partialRound_tempInput_delay_52_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_52_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_52_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_52_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_52_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_52_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_53_valid;
  reg                 partialRound_tempInput_delay_53_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_53_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_53_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_53_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_53_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_53_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_54_valid;
  reg                 partialRound_tempInput_delay_54_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_54_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_54_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_54_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_54_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_54_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_55_valid;
  reg                 partialRound_tempInput_delay_55_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_55_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_55_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_55_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_55_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_55_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_56_valid;
  reg                 partialRound_tempInput_delay_56_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_56_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_56_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_56_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_56_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_56_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_57_valid;
  reg                 partialRound_tempInput_delay_57_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_57_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_57_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_57_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_57_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_57_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_58_valid;
  reg                 partialRound_tempInput_delay_58_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_58_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_58_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_58_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_58_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_58_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_59_valid;
  reg                 partialRound_tempInput_delay_59_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_59_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_59_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_59_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_59_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_59_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_60_valid;
  reg                 partialRound_tempInput_delay_60_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_60_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_60_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_60_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_60_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_60_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_61_valid;
  reg                 partialRound_tempInput_delay_61_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_61_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_61_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_61_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_61_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_61_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_62_valid;
  reg                 partialRound_tempInput_delay_62_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_62_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_62_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_62_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_62_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_62_payload_stateElements_11;
  reg                 partialRound_tempInput_delay_63_valid;
  reg                 partialRound_tempInput_delay_63_payload_isFull;
  reg        [2:0]    partialRound_tempInput_delay_63_payload_fullRound;
  reg        [5:0]    partialRound_tempInput_delay_63_payload_partialRound;
  reg        [3:0]    partialRound_tempInput_delay_63_payload_stateSize;
  reg        [7:0]    partialRound_tempInput_delay_63_payload_stateID;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_0;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_1;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_2;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_3;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_4;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_5;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_6;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_7;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_8;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_9;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_10;
  reg        [254:0]  partialRound_tempInput_delay_63_payload_stateElements_11;
  reg                 partialRound_contextDelayed_valid;
  reg                 partialRound_contextDelayed_payload_isFull;
  reg        [2:0]    partialRound_contextDelayed_payload_fullRound;
  reg        [5:0]    partialRound_contextDelayed_payload_partialRound;
  reg        [3:0]    partialRound_contextDelayed_payload_stateSize;
  reg        [7:0]    partialRound_contextDelayed_payload_stateID;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_0;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_1;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_2;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_3;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_4;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_5;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_6;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_7;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_8;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_9;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_10;
  reg        [254:0]  partialRound_contextDelayed_payload_stateElements_11;
  reg        [254:0]  _zz_partialRound_output_payload_stateElements_0;
  reg        [254:0]  _zz_partialRound_output_payload_stateElements_3;
  reg        [254:0]  _zz_partialRound_output_payload_stateElements_4;
  reg        [254:0]  _zz_partialRound_output_payload_stateElements_5;
  reg        [254:0]  _zz_partialRound_output_payload_stateElements_6;
  reg        [254:0]  _zz_partialRound_output_payload_stateElements_7;
  reg        [254:0]  _zz_partialRound_output_payload_stateElements_8;
  wire                when_MDSMatrixAdders_l91;
  wire                when_MDSMatrixAdders_l94;
  reg                 partialRound_output_valid;
  reg                 partialRound_output_payload_isFull;
  reg        [2:0]    partialRound_output_payload_fullRound;
  reg        [5:0]    partialRound_output_payload_partialRound;
  reg        [3:0]    partialRound_output_payload_stateSize;
  reg        [7:0]    partialRound_output_payload_stateID;
  reg        [254:0]  partialRound_output_payload_stateElements_0;
  reg        [254:0]  partialRound_output_payload_stateElements_1;
  reg        [254:0]  partialRound_output_payload_stateElements_2;
  reg        [254:0]  partialRound_output_payload_stateElements_3;
  reg        [254:0]  partialRound_output_payload_stateElements_4;
  reg        [254:0]  partialRound_output_payload_stateElements_5;
  reg        [254:0]  partialRound_output_payload_stateElements_6;
  reg        [254:0]  partialRound_output_payload_stateElements_7;
  reg        [254:0]  partialRound_output_payload_stateElements_8;
  reg        [254:0]  partialRound_output_payload_stateElements_9;
  reg        [254:0]  partialRound_output_payload_stateElements_10;
  reg        [254:0]  partialRound_output_payload_stateElements_11;
  wire                fullRound_input_valid;
  wire                fullRound_input_payload_isFull;
  wire       [2:0]    fullRound_input_payload_fullRound;
  wire       [5:0]    fullRound_input_payload_partialRound;
  wire       [3:0]    fullRound_input_payload_stateSize;
  wire       [7:0]    fullRound_input_payload_stateID;
  wire       [254:0]  fullRound_input_payload_stateElements_0;
  wire       [254:0]  fullRound_input_payload_stateElements_1;
  wire       [254:0]  fullRound_input_payload_stateElements_2;
  wire       [254:0]  fullRound_input_payload_stateElements_3;
  wire       [254:0]  fullRound_input_payload_stateElements_4;
  wire       [254:0]  fullRound_input_payload_stateElements_5;
  wire       [254:0]  fullRound_input_payload_stateElements_6;
  wire       [254:0]  fullRound_input_payload_stateElements_7;
  wire       [254:0]  fullRound_input_payload_stateElements_8;
  wire       [254:0]  fullRound_input_payload_stateElements_9;
  wire       [254:0]  fullRound_input_payload_stateElements_10;
  wire       [254:0]  fullRound_input_payload_stateElements_11;
  reg                 fullRound_output_valid;
  wire                fullRound_output_payload_isFull;
  wire       [2:0]    fullRound_output_payload_fullRound;
  wire       [5:0]    fullRound_output_payload_partialRound;
  wire       [3:0]    fullRound_output_payload_stateSize;
  wire       [7:0]    fullRound_output_payload_stateID;
  wire       [254:0]  fullRound_output_payload_stateElements_0;
  wire       [254:0]  fullRound_output_payload_stateElements_1;
  wire       [254:0]  fullRound_output_payload_stateElements_2;
  wire       [254:0]  fullRound_output_payload_stateElements_3;
  wire       [254:0]  fullRound_output_payload_stateElements_4;
  wire       [254:0]  fullRound_output_payload_stateElements_5;
  wire       [254:0]  fullRound_output_payload_stateElements_6;
  wire       [254:0]  fullRound_output_payload_stateElements_7;
  wire       [254:0]  fullRound_output_payload_stateElements_8;
  wire       [254:0]  fullRound_output_payload_stateElements_9;
  wire       [254:0]  fullRound_output_payload_stateElements_10;
  wire       [254:0]  fullRound_output_payload_stateElements_11;
  wire                fullRound_adderTreeInput_valid;
  wire       [254:0]  fullRound_adderTreeInput_payload_0;
  wire       [254:0]  fullRound_adderTreeInput_payload_1;
  wire       [254:0]  fullRound_adderTreeInput_payload_2;
  wire       [254:0]  fullRound_adderTreeInput_payload_3;
  wire       [254:0]  fullRound_adderTreeInput_payload_4;
  wire       [254:0]  fullRound_adderTreeInput_payload_5;
  wire       [254:0]  fullRound_adderTreeInput_payload_6;
  wire       [254:0]  fullRound_adderTreeInput_payload_7;
  wire       [254:0]  fullRound_adderTreeInput_payload_8;
  wire       [254:0]  fullRound_adderTreeInput_payload_9;
  wire       [254:0]  fullRound_adderTreeInput_payload_10;
  wire       [254:0]  fullRound_adderTreeInput_payload_11;
  wire                fullRound_addContext_valid;
  wire                fullRound_addContext_payload_isFull;
  wire       [2:0]    fullRound_addContext_payload_fullRound;
  wire       [5:0]    fullRound_addContext_payload_partialRound;
  wire       [3:0]    fullRound_addContext_payload_stateSize;
  wire       [7:0]    fullRound_addContext_payload_stateID;
  reg                 fullRound_addContext_delay_1_valid;
  reg                 fullRound_addContext_delay_1_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_1_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_1_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_1_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_1_payload_stateID;
  reg                 fullRound_addContext_delay_2_valid;
  reg                 fullRound_addContext_delay_2_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_2_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_2_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_2_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_2_payload_stateID;
  reg                 fullRound_addContext_delay_3_valid;
  reg                 fullRound_addContext_delay_3_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_3_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_3_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_3_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_3_payload_stateID;
  reg                 fullRound_addContext_delay_4_valid;
  reg                 fullRound_addContext_delay_4_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_4_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_4_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_4_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_4_payload_stateID;
  reg                 fullRound_addContext_delay_5_valid;
  reg                 fullRound_addContext_delay_5_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_5_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_5_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_5_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_5_payload_stateID;
  reg                 fullRound_addContext_delay_6_valid;
  reg                 fullRound_addContext_delay_6_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_6_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_6_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_6_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_6_payload_stateID;
  reg                 fullRound_addContext_delay_7_valid;
  reg                 fullRound_addContext_delay_7_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_7_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_7_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_7_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_7_payload_stateID;
  reg                 fullRound_addContext_delay_8_valid;
  reg                 fullRound_addContext_delay_8_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_8_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_8_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_8_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_8_payload_stateID;
  reg                 fullRound_addContext_delay_9_valid;
  reg                 fullRound_addContext_delay_9_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_9_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_9_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_9_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_9_payload_stateID;
  reg                 fullRound_addContext_delay_10_valid;
  reg                 fullRound_addContext_delay_10_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_10_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_10_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_10_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_10_payload_stateID;
  reg                 fullRound_addContext_delay_11_valid;
  reg                 fullRound_addContext_delay_11_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_11_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_11_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_11_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_11_payload_stateID;
  reg                 fullRound_addContext_delay_12_valid;
  reg                 fullRound_addContext_delay_12_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_12_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_12_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_12_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_12_payload_stateID;
  reg                 fullRound_addContext_delay_13_valid;
  reg                 fullRound_addContext_delay_13_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_13_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_13_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_13_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_13_payload_stateID;
  reg                 fullRound_addContext_delay_14_valid;
  reg                 fullRound_addContext_delay_14_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_14_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_14_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_14_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_14_payload_stateID;
  reg                 fullRound_addContext_delay_15_valid;
  reg                 fullRound_addContext_delay_15_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_15_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_15_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_15_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_15_payload_stateID;
  reg                 fullRound_addContext_delay_16_valid;
  reg                 fullRound_addContext_delay_16_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_16_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_16_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_16_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_16_payload_stateID;
  reg                 fullRound_addContext_delay_17_valid;
  reg                 fullRound_addContext_delay_17_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_17_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_17_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_17_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_17_payload_stateID;
  reg                 fullRound_addContext_delay_18_valid;
  reg                 fullRound_addContext_delay_18_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_18_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_18_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_18_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_18_payload_stateID;
  reg                 fullRound_addContext_delay_19_valid;
  reg                 fullRound_addContext_delay_19_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_19_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_19_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_19_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_19_payload_stateID;
  reg                 fullRound_addContext_delay_20_valid;
  reg                 fullRound_addContext_delay_20_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_20_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_20_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_20_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_20_payload_stateID;
  reg                 fullRound_addContext_delay_21_valid;
  reg                 fullRound_addContext_delay_21_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_21_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_21_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_21_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_21_payload_stateID;
  reg                 fullRound_addContext_delay_22_valid;
  reg                 fullRound_addContext_delay_22_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_22_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_22_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_22_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_22_payload_stateID;
  reg                 fullRound_addContext_delay_23_valid;
  reg                 fullRound_addContext_delay_23_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_23_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_23_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_23_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_23_payload_stateID;
  reg                 fullRound_addContext_delay_24_valid;
  reg                 fullRound_addContext_delay_24_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_24_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_24_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_24_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_24_payload_stateID;
  reg                 fullRound_addContext_delay_25_valid;
  reg                 fullRound_addContext_delay_25_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_25_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_25_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_25_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_25_payload_stateID;
  reg                 fullRound_addContext_delay_26_valid;
  reg                 fullRound_addContext_delay_26_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_26_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_26_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_26_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_26_payload_stateID;
  reg                 fullRound_addContext_delay_27_valid;
  reg                 fullRound_addContext_delay_27_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_27_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_27_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_27_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_27_payload_stateID;
  reg                 fullRound_addContext_delay_28_valid;
  reg                 fullRound_addContext_delay_28_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_28_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_28_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_28_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_28_payload_stateID;
  reg                 fullRound_addContext_delay_29_valid;
  reg                 fullRound_addContext_delay_29_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_29_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_29_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_29_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_29_payload_stateID;
  reg                 fullRound_addContext_delay_30_valid;
  reg                 fullRound_addContext_delay_30_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_30_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_30_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_30_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_30_payload_stateID;
  reg                 fullRound_addContext_delay_31_valid;
  reg                 fullRound_addContext_delay_31_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_31_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_31_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_31_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_31_payload_stateID;
  reg                 fullRound_addContext_delay_32_valid;
  reg                 fullRound_addContext_delay_32_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_32_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_32_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_32_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_32_payload_stateID;
  reg                 fullRound_addContext_delay_33_valid;
  reg                 fullRound_addContext_delay_33_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_33_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_33_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_33_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_33_payload_stateID;
  reg                 fullRound_addContext_delay_34_valid;
  reg                 fullRound_addContext_delay_34_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_34_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_34_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_34_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_34_payload_stateID;
  reg                 fullRound_addContext_delay_35_valid;
  reg                 fullRound_addContext_delay_35_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_35_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_35_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_35_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_35_payload_stateID;
  reg                 fullRound_addContext_delay_36_valid;
  reg                 fullRound_addContext_delay_36_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_36_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_36_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_36_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_36_payload_stateID;
  reg                 fullRound_addContext_delay_37_valid;
  reg                 fullRound_addContext_delay_37_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_37_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_37_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_37_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_37_payload_stateID;
  reg                 fullRound_addContext_delay_38_valid;
  reg                 fullRound_addContext_delay_38_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_38_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_38_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_38_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_38_payload_stateID;
  reg                 fullRound_addContext_delay_39_valid;
  reg                 fullRound_addContext_delay_39_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_39_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_39_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_39_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_39_payload_stateID;
  reg                 fullRound_addContext_delay_40_valid;
  reg                 fullRound_addContext_delay_40_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_40_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_40_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_40_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_40_payload_stateID;
  reg                 fullRound_addContext_delay_41_valid;
  reg                 fullRound_addContext_delay_41_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_41_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_41_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_41_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_41_payload_stateID;
  reg                 fullRound_addContext_delay_42_valid;
  reg                 fullRound_addContext_delay_42_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_42_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_42_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_42_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_42_payload_stateID;
  reg                 fullRound_addContext_delay_43_valid;
  reg                 fullRound_addContext_delay_43_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_43_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_43_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_43_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_43_payload_stateID;
  reg                 fullRound_addContext_delay_44_valid;
  reg                 fullRound_addContext_delay_44_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_44_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_44_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_44_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_44_payload_stateID;
  reg                 fullRound_addContext_delay_45_valid;
  reg                 fullRound_addContext_delay_45_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_45_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_45_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_45_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_45_payload_stateID;
  reg                 fullRound_addContext_delay_46_valid;
  reg                 fullRound_addContext_delay_46_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_46_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_46_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_46_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_46_payload_stateID;
  reg                 fullRound_addContext_delay_47_valid;
  reg                 fullRound_addContext_delay_47_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_47_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_47_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_47_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_47_payload_stateID;
  reg                 fullRound_addContext_delay_48_valid;
  reg                 fullRound_addContext_delay_48_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_48_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_48_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_48_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_48_payload_stateID;
  reg                 fullRound_addContext_delay_49_valid;
  reg                 fullRound_addContext_delay_49_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_49_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_49_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_49_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_49_payload_stateID;
  reg                 fullRound_addContext_delay_50_valid;
  reg                 fullRound_addContext_delay_50_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_50_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_50_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_50_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_50_payload_stateID;
  reg                 fullRound_addContext_delay_51_valid;
  reg                 fullRound_addContext_delay_51_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_51_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_51_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_51_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_51_payload_stateID;
  reg                 fullRound_addContext_delay_52_valid;
  reg                 fullRound_addContext_delay_52_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_52_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_52_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_52_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_52_payload_stateID;
  reg                 fullRound_addContext_delay_53_valid;
  reg                 fullRound_addContext_delay_53_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_53_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_53_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_53_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_53_payload_stateID;
  reg                 fullRound_addContext_delay_54_valid;
  reg                 fullRound_addContext_delay_54_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_54_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_54_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_54_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_54_payload_stateID;
  reg                 fullRound_addContext_delay_55_valid;
  reg                 fullRound_addContext_delay_55_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_55_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_55_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_55_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_55_payload_stateID;
  reg                 fullRound_addContext_delay_56_valid;
  reg                 fullRound_addContext_delay_56_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_56_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_56_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_56_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_56_payload_stateID;
  reg                 fullRound_addContext_delay_57_valid;
  reg                 fullRound_addContext_delay_57_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_57_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_57_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_57_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_57_payload_stateID;
  reg                 fullRound_addContext_delay_58_valid;
  reg                 fullRound_addContext_delay_58_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_58_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_58_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_58_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_58_payload_stateID;
  reg                 fullRound_addContext_delay_59_valid;
  reg                 fullRound_addContext_delay_59_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_59_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_59_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_59_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_59_payload_stateID;
  reg                 fullRound_addContext_delay_60_valid;
  reg                 fullRound_addContext_delay_60_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_60_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_60_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_60_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_60_payload_stateID;
  reg                 fullRound_addContext_delay_61_valid;
  reg                 fullRound_addContext_delay_61_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_61_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_61_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_61_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_61_payload_stateID;
  reg                 fullRound_addContext_delay_62_valid;
  reg                 fullRound_addContext_delay_62_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_62_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_62_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_62_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_62_payload_stateID;
  reg                 fullRound_addContext_delay_63_valid;
  reg                 fullRound_addContext_delay_63_payload_isFull;
  reg        [2:0]    fullRound_addContext_delay_63_payload_fullRound;
  reg        [5:0]    fullRound_addContext_delay_63_payload_partialRound;
  reg        [3:0]    fullRound_addContext_delay_63_payload_stateSize;
  reg        [7:0]    fullRound_addContext_delay_63_payload_stateID;
  reg                 fullRound_addContextDelayed_valid;
  reg                 fullRound_addContextDelayed_payload_isFull;
  reg        [2:0]    fullRound_addContextDelayed_payload_fullRound;
  reg        [5:0]    fullRound_addContextDelayed_payload_partialRound;
  reg        [3:0]    fullRound_addContextDelayed_payload_stateSize;
  reg        [7:0]    fullRound_addContextDelayed_payload_stateID;
  wire                fullRound_deserialization_wantExit;
  reg                 fullRound_deserialization_wantStart;
  wire                fullRound_deserialization_wantKill;
  reg        [3:0]    fullRound_deserialization_counter;
  reg                 fullRound_deserialization_tempOutput_isFull;
  reg        [2:0]    fullRound_deserialization_tempOutput_fullRound;
  reg        [5:0]    fullRound_deserialization_tempOutput_partialRound;
  reg        [3:0]    fullRound_deserialization_tempOutput_stateSize;
  reg        [7:0]    fullRound_deserialization_tempOutput_stateID;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_0;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_1;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_2;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_3;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_4;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_5;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_6;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_7;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_8;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_9;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_10;
  reg        [254:0]  fullRound_deserialization_tempOutput_stateElements_11;
  wire                fullRound_deserialization_adderTreeValid;
  reg        [1:0]    fullRound_deserialization_stateReg;
  reg        [1:0]    fullRound_deserialization_stateNext;
  wire       [15:0]   _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire                _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire                _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;
  wire                _zz_13;
  wire                when_MDSMatrixAdders_l147;
  wire                when_StateMachine_l222;
  `ifndef SYNTHESIS
  reg [31:0] fullRound_deserialization_stateReg_string;
  reg [31:0] fullRound_deserialization_stateNext_string;
  `endif


  assign _zz_when_MDSMatrixAdders_l147 = (fullRound_deserialization_counter + 4'b0001);
  AdderTree adderTree_1 (
    .io_input_valid         (adderTree_1_io_input_valid              ), //i
    .io_input_payload_0     (adderTree_1_io_input_payload_0[254:0]   ), //i
    .io_input_payload_1     (adderTree_1_io_input_payload_1[254:0]   ), //i
    .io_input_payload_2     (adderTree_1_io_input_payload_2[254:0]   ), //i
    .io_input_payload_3     (adderTree_1_io_input_payload_3[254:0]   ), //i
    .io_input_payload_4     (adderTree_1_io_input_payload_4[254:0]   ), //i
    .io_input_payload_5     (adderTree_1_io_input_payload_5[254:0]   ), //i
    .io_input_payload_6     (adderTree_1_io_input_payload_6[254:0]   ), //i
    .io_input_payload_7     (adderTree_1_io_input_payload_7[254:0]   ), //i
    .io_input_payload_8     (adderTree_1_io_input_payload_8[254:0]   ), //i
    .io_input_payload_9     (adderTree_1_io_input_payload_9[254:0]   ), //i
    .io_input_payload_10    (adderTree_1_io_input_payload_10[254:0]  ), //i
    .io_input_payload_11    (adderTree_1_io_input_payload_11[254:0]  ), //i
    .io_output_valid        (adderTree_1_io_output_valid             ), //o
    .io_output_payload      (adderTree_1_io_output_payload[254:0]    ), //o
    .clk                    (clk                                     ), //i
    .resetn                 (resetn                                  )  //i
  );
  ShiftMatrix fullRound_shiftMat (
    .io_input_valid                        (fullRound_input_valid                                         ), //i
    .io_input_payload_isFull               (fullRound_input_payload_isFull                                ), //i
    .io_input_payload_fullRound            (fullRound_input_payload_fullRound[2:0]                        ), //i
    .io_input_payload_partialRound         (fullRound_input_payload_partialRound[5:0]                     ), //i
    .io_input_payload_stateSize            (fullRound_input_payload_stateSize[3:0]                        ), //i
    .io_input_payload_stateID              (fullRound_input_payload_stateID[7:0]                          ), //i
    .io_input_payload_stateElements_0      (fullRound_input_payload_stateElements_0[254:0]                ), //i
    .io_input_payload_stateElements_1      (fullRound_input_payload_stateElements_1[254:0]                ), //i
    .io_input_payload_stateElements_2      (fullRound_input_payload_stateElements_2[254:0]                ), //i
    .io_input_payload_stateElements_3      (fullRound_input_payload_stateElements_3[254:0]                ), //i
    .io_input_payload_stateElements_4      (fullRound_input_payload_stateElements_4[254:0]                ), //i
    .io_input_payload_stateElements_5      (fullRound_input_payload_stateElements_5[254:0]                ), //i
    .io_input_payload_stateElements_6      (fullRound_input_payload_stateElements_6[254:0]                ), //i
    .io_input_payload_stateElements_7      (fullRound_input_payload_stateElements_7[254:0]                ), //i
    .io_input_payload_stateElements_8      (fullRound_input_payload_stateElements_8[254:0]                ), //i
    .io_input_payload_stateElements_9      (fullRound_input_payload_stateElements_9[254:0]                ), //i
    .io_input_payload_stateElements_10     (fullRound_input_payload_stateElements_10[254:0]               ), //i
    .io_input_payload_stateElements_11     (fullRound_input_payload_stateElements_11[254:0]               ), //i
    .io_output_valid                       (fullRound_shiftMat_io_output_valid                            ), //o
    .io_output_payload_isFull              (fullRound_shiftMat_io_output_payload_isFull                   ), //o
    .io_output_payload_fullRound           (fullRound_shiftMat_io_output_payload_fullRound[2:0]           ), //o
    .io_output_payload_partialRound        (fullRound_shiftMat_io_output_payload_partialRound[5:0]        ), //o
    .io_output_payload_stateSize           (fullRound_shiftMat_io_output_payload_stateSize[3:0]           ), //o
    .io_output_payload_stateID             (fullRound_shiftMat_io_output_payload_stateID[7:0]             ), //o
    .io_output_payload_stateElements_0     (fullRound_shiftMat_io_output_payload_stateElements_0[254:0]   ), //o
    .io_output_payload_stateElements_1     (fullRound_shiftMat_io_output_payload_stateElements_1[254:0]   ), //o
    .io_output_payload_stateElements_2     (fullRound_shiftMat_io_output_payload_stateElements_2[254:0]   ), //o
    .io_output_payload_stateElements_3     (fullRound_shiftMat_io_output_payload_stateElements_3[254:0]   ), //o
    .io_output_payload_stateElements_4     (fullRound_shiftMat_io_output_payload_stateElements_4[254:0]   ), //o
    .io_output_payload_stateElements_5     (fullRound_shiftMat_io_output_payload_stateElements_5[254:0]   ), //o
    .io_output_payload_stateElements_6     (fullRound_shiftMat_io_output_payload_stateElements_6[254:0]   ), //o
    .io_output_payload_stateElements_7     (fullRound_shiftMat_io_output_payload_stateElements_7[254:0]   ), //o
    .io_output_payload_stateElements_8     (fullRound_shiftMat_io_output_payload_stateElements_8[254:0]   ), //o
    .io_output_payload_stateElements_9     (fullRound_shiftMat_io_output_payload_stateElements_9[254:0]   ), //o
    .io_output_payload_stateElements_10    (fullRound_shiftMat_io_output_payload_stateElements_10[254:0]  ), //o
    .io_output_payload_stateElements_11    (fullRound_shiftMat_io_output_payload_stateElements_11[254:0]  ), //o
    .clk                                   (clk                                                           ), //i
    .resetn                                (resetn                                                        )  //i
  );
  always @(*) begin
    case(_zz_partialRound_bufferOutMuxed_valid_2)
      2'b00 : begin
        _zz_partialRound_bufferOutMuxed_valid_3 = partialRound_bufferOut_0_valid;
        _zz_partialRound_bufferOutMuxed_payload_isFull = partialRound_bufferOut_0_payload_isFull;
        _zz_partialRound_bufferOutMuxed_payload_fullRound = partialRound_bufferOut_0_payload_fullRound;
        _zz_partialRound_bufferOutMuxed_payload_partialRound = partialRound_bufferOut_0_payload_partialRound;
        _zz_partialRound_bufferOutMuxed_payload_stateSize = partialRound_bufferOut_0_payload_stateSize;
        _zz_partialRound_bufferOutMuxed_payload_stateID = partialRound_bufferOut_0_payload_stateID;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_0 = partialRound_bufferOut_0_payload_stateElements_0;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_1 = partialRound_bufferOut_0_payload_stateElements_1;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_2 = partialRound_bufferOut_0_payload_stateElements_2;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_3 = partialRound_bufferOut_0_payload_stateElements_3;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_4 = partialRound_bufferOut_0_payload_stateElements_4;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_5 = partialRound_bufferOut_0_payload_stateElements_5;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_6 = partialRound_bufferOut_0_payload_stateElements_6;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_7 = partialRound_bufferOut_0_payload_stateElements_7;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_8 = partialRound_bufferOut_0_payload_stateElements_8;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_9 = partialRound_bufferOut_0_payload_stateElements_9;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_10 = partialRound_bufferOut_0_payload_stateElements_10;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_11 = partialRound_bufferOut_0_payload_stateElements_11;
      end
      2'b01 : begin
        _zz_partialRound_bufferOutMuxed_valid_3 = partialRound_bufferOut_1_valid;
        _zz_partialRound_bufferOutMuxed_payload_isFull = partialRound_bufferOut_1_payload_isFull;
        _zz_partialRound_bufferOutMuxed_payload_fullRound = partialRound_bufferOut_1_payload_fullRound;
        _zz_partialRound_bufferOutMuxed_payload_partialRound = partialRound_bufferOut_1_payload_partialRound;
        _zz_partialRound_bufferOutMuxed_payload_stateSize = partialRound_bufferOut_1_payload_stateSize;
        _zz_partialRound_bufferOutMuxed_payload_stateID = partialRound_bufferOut_1_payload_stateID;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_0 = partialRound_bufferOut_1_payload_stateElements_0;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_1 = partialRound_bufferOut_1_payload_stateElements_1;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_2 = partialRound_bufferOut_1_payload_stateElements_2;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_3 = partialRound_bufferOut_1_payload_stateElements_3;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_4 = partialRound_bufferOut_1_payload_stateElements_4;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_5 = partialRound_bufferOut_1_payload_stateElements_5;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_6 = partialRound_bufferOut_1_payload_stateElements_6;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_7 = partialRound_bufferOut_1_payload_stateElements_7;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_8 = partialRound_bufferOut_1_payload_stateElements_8;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_9 = partialRound_bufferOut_1_payload_stateElements_9;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_10 = partialRound_bufferOut_1_payload_stateElements_10;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_11 = partialRound_bufferOut_1_payload_stateElements_11;
      end
      2'b10 : begin
        _zz_partialRound_bufferOutMuxed_valid_3 = partialRound_bufferOut_2_valid;
        _zz_partialRound_bufferOutMuxed_payload_isFull = partialRound_bufferOut_2_payload_isFull;
        _zz_partialRound_bufferOutMuxed_payload_fullRound = partialRound_bufferOut_2_payload_fullRound;
        _zz_partialRound_bufferOutMuxed_payload_partialRound = partialRound_bufferOut_2_payload_partialRound;
        _zz_partialRound_bufferOutMuxed_payload_stateSize = partialRound_bufferOut_2_payload_stateSize;
        _zz_partialRound_bufferOutMuxed_payload_stateID = partialRound_bufferOut_2_payload_stateID;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_0 = partialRound_bufferOut_2_payload_stateElements_0;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_1 = partialRound_bufferOut_2_payload_stateElements_1;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_2 = partialRound_bufferOut_2_payload_stateElements_2;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_3 = partialRound_bufferOut_2_payload_stateElements_3;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_4 = partialRound_bufferOut_2_payload_stateElements_4;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_5 = partialRound_bufferOut_2_payload_stateElements_5;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_6 = partialRound_bufferOut_2_payload_stateElements_6;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_7 = partialRound_bufferOut_2_payload_stateElements_7;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_8 = partialRound_bufferOut_2_payload_stateElements_8;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_9 = partialRound_bufferOut_2_payload_stateElements_9;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_10 = partialRound_bufferOut_2_payload_stateElements_10;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_11 = partialRound_bufferOut_2_payload_stateElements_11;
      end
      default : begin
        _zz_partialRound_bufferOutMuxed_valid_3 = partialRound_bufferOut_3_valid;
        _zz_partialRound_bufferOutMuxed_payload_isFull = partialRound_bufferOut_3_payload_isFull;
        _zz_partialRound_bufferOutMuxed_payload_fullRound = partialRound_bufferOut_3_payload_fullRound;
        _zz_partialRound_bufferOutMuxed_payload_partialRound = partialRound_bufferOut_3_payload_partialRound;
        _zz_partialRound_bufferOutMuxed_payload_stateSize = partialRound_bufferOut_3_payload_stateSize;
        _zz_partialRound_bufferOutMuxed_payload_stateID = partialRound_bufferOut_3_payload_stateID;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_0 = partialRound_bufferOut_3_payload_stateElements_0;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_1 = partialRound_bufferOut_3_payload_stateElements_1;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_2 = partialRound_bufferOut_3_payload_stateElements_2;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_3 = partialRound_bufferOut_3_payload_stateElements_3;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_4 = partialRound_bufferOut_3_payload_stateElements_4;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_5 = partialRound_bufferOut_3_payload_stateElements_5;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_6 = partialRound_bufferOut_3_payload_stateElements_6;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_7 = partialRound_bufferOut_3_payload_stateElements_7;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_8 = partialRound_bufferOut_3_payload_stateElements_8;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_9 = partialRound_bufferOut_3_payload_stateElements_9;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_10 = partialRound_bufferOut_3_payload_stateElements_10;
        _zz_partialRound_bufferOutMuxed_payload_stateElements_11 = partialRound_bufferOut_3_payload_stateElements_11;
      end
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(fullRound_deserialization_stateReg)
      fullRound_deserialization_enumDef_BOOT : fullRound_deserialization_stateReg_string = "BOOT";
      fullRound_deserialization_enumDef_IDLE : fullRound_deserialization_stateReg_string = "IDLE";
      fullRound_deserialization_enumDef_BUSY : fullRound_deserialization_stateReg_string = "BUSY";
      fullRound_deserialization_enumDef_DONE : fullRound_deserialization_stateReg_string = "DONE";
      default : fullRound_deserialization_stateReg_string = "????";
    endcase
  end
  always @(*) begin
    case(fullRound_deserialization_stateNext)
      fullRound_deserialization_enumDef_BOOT : fullRound_deserialization_stateNext_string = "BOOT";
      fullRound_deserialization_enumDef_IDLE : fullRound_deserialization_stateNext_string = "IDLE";
      fullRound_deserialization_enumDef_BUSY : fullRound_deserialization_stateNext_string = "BUSY";
      fullRound_deserialization_enumDef_DONE : fullRound_deserialization_stateNext_string = "DONE";
      default : fullRound_deserialization_stateNext_string = "????";
    endcase
  end
  `endif

  assign partialRound_input_valid = (io_input_valid && (! io_input_payload_isFull));
  assign partialRound_input_payload_isFull = io_input_payload_isFull;
  assign partialRound_input_payload_fullRound = io_input_payload_fullRound;
  assign partialRound_input_payload_partialRound = io_input_payload_partialRound;
  assign partialRound_input_payload_stateSize = io_input_payload_stateSize;
  assign partialRound_input_payload_stateID = io_input_payload_stateID;
  assign partialRound_input_payload_stateElements_0 = io_input_payload_stateElements_0;
  assign partialRound_input_payload_stateElements_1 = io_input_payload_stateElements_1;
  assign partialRound_input_payload_stateElements_2 = io_input_payload_stateElements_2;
  assign partialRound_input_payload_stateElements_3 = io_input_payload_stateElements_3;
  assign partialRound_input_payload_stateElements_4 = io_input_payload_stateElements_4;
  assign partialRound_input_payload_stateElements_5 = io_input_payload_stateElements_5;
  assign partialRound_input_payload_stateElements_6 = io_input_payload_stateElements_6;
  assign partialRound_input_payload_stateElements_7 = io_input_payload_stateElements_7;
  assign partialRound_input_payload_stateElements_8 = io_input_payload_stateElements_8;
  assign partialRound_input_payload_stateElements_9 = io_input_payload_stateElements_9;
  assign partialRound_input_payload_stateElements_10 = io_input_payload_stateElements_10;
  assign partialRound_input_payload_stateElements_11 = io_input_payload_stateElements_11;
  assign partialRound_inputBuffered_0_valid = partialRound_input_regNext_valid;
  assign partialRound_inputBuffered_0_payload_isFull = partialRound_input_regNext_payload_isFull;
  assign partialRound_inputBuffered_0_payload_fullRound = partialRound_input_regNext_payload_fullRound;
  assign partialRound_inputBuffered_0_payload_partialRound = partialRound_input_regNext_payload_partialRound;
  assign partialRound_inputBuffered_0_payload_stateSize = partialRound_input_regNext_payload_stateSize;
  assign partialRound_inputBuffered_0_payload_stateID = partialRound_input_regNext_payload_stateID;
  assign partialRound_inputBuffered_0_payload_stateElements_0 = partialRound_input_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_0_payload_stateElements_1 = partialRound_input_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_0_payload_stateElements_2 = partialRound_input_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_0_payload_stateElements_3 = partialRound_input_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_0_payload_stateElements_4 = partialRound_input_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_0_payload_stateElements_5 = partialRound_input_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_0_payload_stateElements_6 = partialRound_input_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_0_payload_stateElements_7 = partialRound_input_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_0_payload_stateElements_8 = partialRound_input_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_0_payload_stateElements_9 = partialRound_input_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_0_payload_stateElements_10 = partialRound_input_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_0_payload_stateElements_11 = partialRound_input_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_1_valid = partialRound_inputBuffered_0_regNext_valid;
  assign partialRound_inputBuffered_1_payload_isFull = partialRound_inputBuffered_0_regNext_payload_isFull;
  assign partialRound_inputBuffered_1_payload_fullRound = partialRound_inputBuffered_0_regNext_payload_fullRound;
  assign partialRound_inputBuffered_1_payload_partialRound = partialRound_inputBuffered_0_regNext_payload_partialRound;
  assign partialRound_inputBuffered_1_payload_stateSize = partialRound_inputBuffered_0_regNext_payload_stateSize;
  assign partialRound_inputBuffered_1_payload_stateID = partialRound_inputBuffered_0_regNext_payload_stateID;
  assign partialRound_inputBuffered_1_payload_stateElements_0 = partialRound_inputBuffered_0_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_1_payload_stateElements_1 = partialRound_inputBuffered_0_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_1_payload_stateElements_2 = partialRound_inputBuffered_0_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_1_payload_stateElements_3 = partialRound_inputBuffered_0_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_1_payload_stateElements_4 = partialRound_inputBuffered_0_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_1_payload_stateElements_5 = partialRound_inputBuffered_0_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_1_payload_stateElements_6 = partialRound_inputBuffered_0_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_1_payload_stateElements_7 = partialRound_inputBuffered_0_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_1_payload_stateElements_8 = partialRound_inputBuffered_0_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_1_payload_stateElements_9 = partialRound_inputBuffered_0_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_1_payload_stateElements_10 = partialRound_inputBuffered_0_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_1_payload_stateElements_11 = partialRound_inputBuffered_0_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_2_valid = partialRound_inputBuffered_1_regNext_valid;
  assign partialRound_inputBuffered_2_payload_isFull = partialRound_inputBuffered_1_regNext_payload_isFull;
  assign partialRound_inputBuffered_2_payload_fullRound = partialRound_inputBuffered_1_regNext_payload_fullRound;
  assign partialRound_inputBuffered_2_payload_partialRound = partialRound_inputBuffered_1_regNext_payload_partialRound;
  assign partialRound_inputBuffered_2_payload_stateSize = partialRound_inputBuffered_1_regNext_payload_stateSize;
  assign partialRound_inputBuffered_2_payload_stateID = partialRound_inputBuffered_1_regNext_payload_stateID;
  assign partialRound_inputBuffered_2_payload_stateElements_0 = partialRound_inputBuffered_1_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_2_payload_stateElements_1 = partialRound_inputBuffered_1_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_2_payload_stateElements_2 = partialRound_inputBuffered_1_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_2_payload_stateElements_3 = partialRound_inputBuffered_1_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_2_payload_stateElements_4 = partialRound_inputBuffered_1_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_2_payload_stateElements_5 = partialRound_inputBuffered_1_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_2_payload_stateElements_6 = partialRound_inputBuffered_1_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_2_payload_stateElements_7 = partialRound_inputBuffered_1_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_2_payload_stateElements_8 = partialRound_inputBuffered_1_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_2_payload_stateElements_9 = partialRound_inputBuffered_1_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_2_payload_stateElements_10 = partialRound_inputBuffered_1_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_2_payload_stateElements_11 = partialRound_inputBuffered_1_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_3_valid = partialRound_inputBuffered_2_regNext_valid;
  assign partialRound_inputBuffered_3_payload_isFull = partialRound_inputBuffered_2_regNext_payload_isFull;
  assign partialRound_inputBuffered_3_payload_fullRound = partialRound_inputBuffered_2_regNext_payload_fullRound;
  assign partialRound_inputBuffered_3_payload_partialRound = partialRound_inputBuffered_2_regNext_payload_partialRound;
  assign partialRound_inputBuffered_3_payload_stateSize = partialRound_inputBuffered_2_regNext_payload_stateSize;
  assign partialRound_inputBuffered_3_payload_stateID = partialRound_inputBuffered_2_regNext_payload_stateID;
  assign partialRound_inputBuffered_3_payload_stateElements_0 = partialRound_inputBuffered_2_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_3_payload_stateElements_1 = partialRound_inputBuffered_2_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_3_payload_stateElements_2 = partialRound_inputBuffered_2_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_3_payload_stateElements_3 = partialRound_inputBuffered_2_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_3_payload_stateElements_4 = partialRound_inputBuffered_2_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_3_payload_stateElements_5 = partialRound_inputBuffered_2_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_3_payload_stateElements_6 = partialRound_inputBuffered_2_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_3_payload_stateElements_7 = partialRound_inputBuffered_2_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_3_payload_stateElements_8 = partialRound_inputBuffered_2_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_3_payload_stateElements_9 = partialRound_inputBuffered_2_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_3_payload_stateElements_10 = partialRound_inputBuffered_2_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_3_payload_stateElements_11 = partialRound_inputBuffered_2_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_4_valid = partialRound_inputBuffered_3_regNext_valid;
  assign partialRound_inputBuffered_4_payload_isFull = partialRound_inputBuffered_3_regNext_payload_isFull;
  assign partialRound_inputBuffered_4_payload_fullRound = partialRound_inputBuffered_3_regNext_payload_fullRound;
  assign partialRound_inputBuffered_4_payload_partialRound = partialRound_inputBuffered_3_regNext_payload_partialRound;
  assign partialRound_inputBuffered_4_payload_stateSize = partialRound_inputBuffered_3_regNext_payload_stateSize;
  assign partialRound_inputBuffered_4_payload_stateID = partialRound_inputBuffered_3_regNext_payload_stateID;
  assign partialRound_inputBuffered_4_payload_stateElements_0 = partialRound_inputBuffered_3_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_4_payload_stateElements_1 = partialRound_inputBuffered_3_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_4_payload_stateElements_2 = partialRound_inputBuffered_3_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_4_payload_stateElements_3 = partialRound_inputBuffered_3_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_4_payload_stateElements_4 = partialRound_inputBuffered_3_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_4_payload_stateElements_5 = partialRound_inputBuffered_3_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_4_payload_stateElements_6 = partialRound_inputBuffered_3_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_4_payload_stateElements_7 = partialRound_inputBuffered_3_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_4_payload_stateElements_8 = partialRound_inputBuffered_3_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_4_payload_stateElements_9 = partialRound_inputBuffered_3_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_4_payload_stateElements_10 = partialRound_inputBuffered_3_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_4_payload_stateElements_11 = partialRound_inputBuffered_3_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_5_valid = partialRound_inputBuffered_4_regNext_valid;
  assign partialRound_inputBuffered_5_payload_isFull = partialRound_inputBuffered_4_regNext_payload_isFull;
  assign partialRound_inputBuffered_5_payload_fullRound = partialRound_inputBuffered_4_regNext_payload_fullRound;
  assign partialRound_inputBuffered_5_payload_partialRound = partialRound_inputBuffered_4_regNext_payload_partialRound;
  assign partialRound_inputBuffered_5_payload_stateSize = partialRound_inputBuffered_4_regNext_payload_stateSize;
  assign partialRound_inputBuffered_5_payload_stateID = partialRound_inputBuffered_4_regNext_payload_stateID;
  assign partialRound_inputBuffered_5_payload_stateElements_0 = partialRound_inputBuffered_4_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_5_payload_stateElements_1 = partialRound_inputBuffered_4_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_5_payload_stateElements_2 = partialRound_inputBuffered_4_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_5_payload_stateElements_3 = partialRound_inputBuffered_4_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_5_payload_stateElements_4 = partialRound_inputBuffered_4_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_5_payload_stateElements_5 = partialRound_inputBuffered_4_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_5_payload_stateElements_6 = partialRound_inputBuffered_4_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_5_payload_stateElements_7 = partialRound_inputBuffered_4_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_5_payload_stateElements_8 = partialRound_inputBuffered_4_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_5_payload_stateElements_9 = partialRound_inputBuffered_4_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_5_payload_stateElements_10 = partialRound_inputBuffered_4_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_5_payload_stateElements_11 = partialRound_inputBuffered_4_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_6_valid = partialRound_inputBuffered_5_regNext_valid;
  assign partialRound_inputBuffered_6_payload_isFull = partialRound_inputBuffered_5_regNext_payload_isFull;
  assign partialRound_inputBuffered_6_payload_fullRound = partialRound_inputBuffered_5_regNext_payload_fullRound;
  assign partialRound_inputBuffered_6_payload_partialRound = partialRound_inputBuffered_5_regNext_payload_partialRound;
  assign partialRound_inputBuffered_6_payload_stateSize = partialRound_inputBuffered_5_regNext_payload_stateSize;
  assign partialRound_inputBuffered_6_payload_stateID = partialRound_inputBuffered_5_regNext_payload_stateID;
  assign partialRound_inputBuffered_6_payload_stateElements_0 = partialRound_inputBuffered_5_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_6_payload_stateElements_1 = partialRound_inputBuffered_5_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_6_payload_stateElements_2 = partialRound_inputBuffered_5_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_6_payload_stateElements_3 = partialRound_inputBuffered_5_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_6_payload_stateElements_4 = partialRound_inputBuffered_5_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_6_payload_stateElements_5 = partialRound_inputBuffered_5_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_6_payload_stateElements_6 = partialRound_inputBuffered_5_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_6_payload_stateElements_7 = partialRound_inputBuffered_5_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_6_payload_stateElements_8 = partialRound_inputBuffered_5_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_6_payload_stateElements_9 = partialRound_inputBuffered_5_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_6_payload_stateElements_10 = partialRound_inputBuffered_5_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_6_payload_stateElements_11 = partialRound_inputBuffered_5_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_7_valid = partialRound_inputBuffered_6_regNext_valid;
  assign partialRound_inputBuffered_7_payload_isFull = partialRound_inputBuffered_6_regNext_payload_isFull;
  assign partialRound_inputBuffered_7_payload_fullRound = partialRound_inputBuffered_6_regNext_payload_fullRound;
  assign partialRound_inputBuffered_7_payload_partialRound = partialRound_inputBuffered_6_regNext_payload_partialRound;
  assign partialRound_inputBuffered_7_payload_stateSize = partialRound_inputBuffered_6_regNext_payload_stateSize;
  assign partialRound_inputBuffered_7_payload_stateID = partialRound_inputBuffered_6_regNext_payload_stateID;
  assign partialRound_inputBuffered_7_payload_stateElements_0 = partialRound_inputBuffered_6_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_7_payload_stateElements_1 = partialRound_inputBuffered_6_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_7_payload_stateElements_2 = partialRound_inputBuffered_6_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_7_payload_stateElements_3 = partialRound_inputBuffered_6_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_7_payload_stateElements_4 = partialRound_inputBuffered_6_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_7_payload_stateElements_5 = partialRound_inputBuffered_6_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_7_payload_stateElements_6 = partialRound_inputBuffered_6_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_7_payload_stateElements_7 = partialRound_inputBuffered_6_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_7_payload_stateElements_8 = partialRound_inputBuffered_6_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_7_payload_stateElements_9 = partialRound_inputBuffered_6_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_7_payload_stateElements_10 = partialRound_inputBuffered_6_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_7_payload_stateElements_11 = partialRound_inputBuffered_6_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_8_valid = partialRound_inputBuffered_7_regNext_valid;
  assign partialRound_inputBuffered_8_payload_isFull = partialRound_inputBuffered_7_regNext_payload_isFull;
  assign partialRound_inputBuffered_8_payload_fullRound = partialRound_inputBuffered_7_regNext_payload_fullRound;
  assign partialRound_inputBuffered_8_payload_partialRound = partialRound_inputBuffered_7_regNext_payload_partialRound;
  assign partialRound_inputBuffered_8_payload_stateSize = partialRound_inputBuffered_7_regNext_payload_stateSize;
  assign partialRound_inputBuffered_8_payload_stateID = partialRound_inputBuffered_7_regNext_payload_stateID;
  assign partialRound_inputBuffered_8_payload_stateElements_0 = partialRound_inputBuffered_7_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_8_payload_stateElements_1 = partialRound_inputBuffered_7_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_8_payload_stateElements_2 = partialRound_inputBuffered_7_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_8_payload_stateElements_3 = partialRound_inputBuffered_7_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_8_payload_stateElements_4 = partialRound_inputBuffered_7_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_8_payload_stateElements_5 = partialRound_inputBuffered_7_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_8_payload_stateElements_6 = partialRound_inputBuffered_7_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_8_payload_stateElements_7 = partialRound_inputBuffered_7_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_8_payload_stateElements_8 = partialRound_inputBuffered_7_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_8_payload_stateElements_9 = partialRound_inputBuffered_7_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_8_payload_stateElements_10 = partialRound_inputBuffered_7_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_8_payload_stateElements_11 = partialRound_inputBuffered_7_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_9_valid = partialRound_inputBuffered_8_regNext_valid;
  assign partialRound_inputBuffered_9_payload_isFull = partialRound_inputBuffered_8_regNext_payload_isFull;
  assign partialRound_inputBuffered_9_payload_fullRound = partialRound_inputBuffered_8_regNext_payload_fullRound;
  assign partialRound_inputBuffered_9_payload_partialRound = partialRound_inputBuffered_8_regNext_payload_partialRound;
  assign partialRound_inputBuffered_9_payload_stateSize = partialRound_inputBuffered_8_regNext_payload_stateSize;
  assign partialRound_inputBuffered_9_payload_stateID = partialRound_inputBuffered_8_regNext_payload_stateID;
  assign partialRound_inputBuffered_9_payload_stateElements_0 = partialRound_inputBuffered_8_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_9_payload_stateElements_1 = partialRound_inputBuffered_8_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_9_payload_stateElements_2 = partialRound_inputBuffered_8_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_9_payload_stateElements_3 = partialRound_inputBuffered_8_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_9_payload_stateElements_4 = partialRound_inputBuffered_8_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_9_payload_stateElements_5 = partialRound_inputBuffered_8_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_9_payload_stateElements_6 = partialRound_inputBuffered_8_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_9_payload_stateElements_7 = partialRound_inputBuffered_8_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_9_payload_stateElements_8 = partialRound_inputBuffered_8_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_9_payload_stateElements_9 = partialRound_inputBuffered_8_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_9_payload_stateElements_10 = partialRound_inputBuffered_8_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_9_payload_stateElements_11 = partialRound_inputBuffered_8_regNext_payload_stateElements_11;
  assign partialRound_inputBuffered_10_valid = partialRound_inputBuffered_9_regNext_valid;
  assign partialRound_inputBuffered_10_payload_isFull = partialRound_inputBuffered_9_regNext_payload_isFull;
  assign partialRound_inputBuffered_10_payload_fullRound = partialRound_inputBuffered_9_regNext_payload_fullRound;
  assign partialRound_inputBuffered_10_payload_partialRound = partialRound_inputBuffered_9_regNext_payload_partialRound;
  assign partialRound_inputBuffered_10_payload_stateSize = partialRound_inputBuffered_9_regNext_payload_stateSize;
  assign partialRound_inputBuffered_10_payload_stateID = partialRound_inputBuffered_9_regNext_payload_stateID;
  assign partialRound_inputBuffered_10_payload_stateElements_0 = partialRound_inputBuffered_9_regNext_payload_stateElements_0;
  assign partialRound_inputBuffered_10_payload_stateElements_1 = partialRound_inputBuffered_9_regNext_payload_stateElements_1;
  assign partialRound_inputBuffered_10_payload_stateElements_2 = partialRound_inputBuffered_9_regNext_payload_stateElements_2;
  assign partialRound_inputBuffered_10_payload_stateElements_3 = partialRound_inputBuffered_9_regNext_payload_stateElements_3;
  assign partialRound_inputBuffered_10_payload_stateElements_4 = partialRound_inputBuffered_9_regNext_payload_stateElements_4;
  assign partialRound_inputBuffered_10_payload_stateElements_5 = partialRound_inputBuffered_9_regNext_payload_stateElements_5;
  assign partialRound_inputBuffered_10_payload_stateElements_6 = partialRound_inputBuffered_9_regNext_payload_stateElements_6;
  assign partialRound_inputBuffered_10_payload_stateElements_7 = partialRound_inputBuffered_9_regNext_payload_stateElements_7;
  assign partialRound_inputBuffered_10_payload_stateElements_8 = partialRound_inputBuffered_9_regNext_payload_stateElements_8;
  assign partialRound_inputBuffered_10_payload_stateElements_9 = partialRound_inputBuffered_9_regNext_payload_stateElements_9;
  assign partialRound_inputBuffered_10_payload_stateElements_10 = partialRound_inputBuffered_9_regNext_payload_stateElements_10;
  assign partialRound_inputBuffered_10_payload_stateElements_11 = partialRound_inputBuffered_9_regNext_payload_stateElements_11;
  assign partialRound_bufferOut_0_valid = (partialRound_inputBuffered_1_valid && (partialRound_inputBuffered_1_payload_stateSize == 4'b0011));
  assign partialRound_bufferOut_0_payload_isFull = partialRound_inputBuffered_1_payload_isFull;
  assign partialRound_bufferOut_0_payload_fullRound = partialRound_inputBuffered_1_payload_fullRound;
  assign partialRound_bufferOut_0_payload_partialRound = partialRound_inputBuffered_1_payload_partialRound;
  assign partialRound_bufferOut_0_payload_stateSize = partialRound_inputBuffered_1_payload_stateSize;
  assign partialRound_bufferOut_0_payload_stateID = partialRound_inputBuffered_1_payload_stateID;
  assign partialRound_bufferOut_0_payload_stateElements_0 = partialRound_inputBuffered_1_payload_stateElements_0;
  assign partialRound_bufferOut_0_payload_stateElements_1 = partialRound_inputBuffered_1_payload_stateElements_1;
  assign partialRound_bufferOut_0_payload_stateElements_2 = partialRound_inputBuffered_1_payload_stateElements_2;
  assign partialRound_bufferOut_0_payload_stateElements_3 = partialRound_inputBuffered_1_payload_stateElements_3;
  assign partialRound_bufferOut_0_payload_stateElements_4 = partialRound_inputBuffered_1_payload_stateElements_4;
  assign partialRound_bufferOut_0_payload_stateElements_5 = partialRound_inputBuffered_1_payload_stateElements_5;
  assign partialRound_bufferOut_0_payload_stateElements_6 = partialRound_inputBuffered_1_payload_stateElements_6;
  assign partialRound_bufferOut_0_payload_stateElements_7 = partialRound_inputBuffered_1_payload_stateElements_7;
  assign partialRound_bufferOut_0_payload_stateElements_8 = partialRound_inputBuffered_1_payload_stateElements_8;
  assign partialRound_bufferOut_0_payload_stateElements_9 = partialRound_inputBuffered_1_payload_stateElements_9;
  assign partialRound_bufferOut_0_payload_stateElements_10 = partialRound_inputBuffered_1_payload_stateElements_10;
  assign partialRound_bufferOut_0_payload_stateElements_11 = partialRound_inputBuffered_1_payload_stateElements_11;
  assign partialRound_bufferOut_1_valid = (partialRound_inputBuffered_3_valid && (partialRound_inputBuffered_3_payload_stateSize == 4'b0101));
  assign partialRound_bufferOut_1_payload_isFull = partialRound_inputBuffered_3_payload_isFull;
  assign partialRound_bufferOut_1_payload_fullRound = partialRound_inputBuffered_3_payload_fullRound;
  assign partialRound_bufferOut_1_payload_partialRound = partialRound_inputBuffered_3_payload_partialRound;
  assign partialRound_bufferOut_1_payload_stateSize = partialRound_inputBuffered_3_payload_stateSize;
  assign partialRound_bufferOut_1_payload_stateID = partialRound_inputBuffered_3_payload_stateID;
  assign partialRound_bufferOut_1_payload_stateElements_0 = partialRound_inputBuffered_3_payload_stateElements_0;
  assign partialRound_bufferOut_1_payload_stateElements_1 = partialRound_inputBuffered_3_payload_stateElements_1;
  assign partialRound_bufferOut_1_payload_stateElements_2 = partialRound_inputBuffered_3_payload_stateElements_2;
  assign partialRound_bufferOut_1_payload_stateElements_3 = partialRound_inputBuffered_3_payload_stateElements_3;
  assign partialRound_bufferOut_1_payload_stateElements_4 = partialRound_inputBuffered_3_payload_stateElements_4;
  assign partialRound_bufferOut_1_payload_stateElements_5 = partialRound_inputBuffered_3_payload_stateElements_5;
  assign partialRound_bufferOut_1_payload_stateElements_6 = partialRound_inputBuffered_3_payload_stateElements_6;
  assign partialRound_bufferOut_1_payload_stateElements_7 = partialRound_inputBuffered_3_payload_stateElements_7;
  assign partialRound_bufferOut_1_payload_stateElements_8 = partialRound_inputBuffered_3_payload_stateElements_8;
  assign partialRound_bufferOut_1_payload_stateElements_9 = partialRound_inputBuffered_3_payload_stateElements_9;
  assign partialRound_bufferOut_1_payload_stateElements_10 = partialRound_inputBuffered_3_payload_stateElements_10;
  assign partialRound_bufferOut_1_payload_stateElements_11 = partialRound_inputBuffered_3_payload_stateElements_11;
  assign partialRound_bufferOut_2_valid = (partialRound_inputBuffered_7_valid && (partialRound_inputBuffered_7_payload_stateSize == 4'b1001));
  assign partialRound_bufferOut_2_payload_isFull = partialRound_inputBuffered_7_payload_isFull;
  assign partialRound_bufferOut_2_payload_fullRound = partialRound_inputBuffered_7_payload_fullRound;
  assign partialRound_bufferOut_2_payload_partialRound = partialRound_inputBuffered_7_payload_partialRound;
  assign partialRound_bufferOut_2_payload_stateSize = partialRound_inputBuffered_7_payload_stateSize;
  assign partialRound_bufferOut_2_payload_stateID = partialRound_inputBuffered_7_payload_stateID;
  assign partialRound_bufferOut_2_payload_stateElements_0 = partialRound_inputBuffered_7_payload_stateElements_0;
  assign partialRound_bufferOut_2_payload_stateElements_1 = partialRound_inputBuffered_7_payload_stateElements_1;
  assign partialRound_bufferOut_2_payload_stateElements_2 = partialRound_inputBuffered_7_payload_stateElements_2;
  assign partialRound_bufferOut_2_payload_stateElements_3 = partialRound_inputBuffered_7_payload_stateElements_3;
  assign partialRound_bufferOut_2_payload_stateElements_4 = partialRound_inputBuffered_7_payload_stateElements_4;
  assign partialRound_bufferOut_2_payload_stateElements_5 = partialRound_inputBuffered_7_payload_stateElements_5;
  assign partialRound_bufferOut_2_payload_stateElements_6 = partialRound_inputBuffered_7_payload_stateElements_6;
  assign partialRound_bufferOut_2_payload_stateElements_7 = partialRound_inputBuffered_7_payload_stateElements_7;
  assign partialRound_bufferOut_2_payload_stateElements_8 = partialRound_inputBuffered_7_payload_stateElements_8;
  assign partialRound_bufferOut_2_payload_stateElements_9 = partialRound_inputBuffered_7_payload_stateElements_9;
  assign partialRound_bufferOut_2_payload_stateElements_10 = partialRound_inputBuffered_7_payload_stateElements_10;
  assign partialRound_bufferOut_2_payload_stateElements_11 = partialRound_inputBuffered_7_payload_stateElements_11;
  assign partialRound_bufferOut_3_valid = (partialRound_inputBuffered_10_valid && (partialRound_inputBuffered_10_payload_stateSize == 4'b1100));
  assign partialRound_bufferOut_3_payload_isFull = partialRound_inputBuffered_10_payload_isFull;
  assign partialRound_bufferOut_3_payload_fullRound = partialRound_inputBuffered_10_payload_fullRound;
  assign partialRound_bufferOut_3_payload_partialRound = partialRound_inputBuffered_10_payload_partialRound;
  assign partialRound_bufferOut_3_payload_stateSize = partialRound_inputBuffered_10_payload_stateSize;
  assign partialRound_bufferOut_3_payload_stateID = partialRound_inputBuffered_10_payload_stateID;
  assign partialRound_bufferOut_3_payload_stateElements_0 = partialRound_inputBuffered_10_payload_stateElements_0;
  assign partialRound_bufferOut_3_payload_stateElements_1 = partialRound_inputBuffered_10_payload_stateElements_1;
  assign partialRound_bufferOut_3_payload_stateElements_2 = partialRound_inputBuffered_10_payload_stateElements_2;
  assign partialRound_bufferOut_3_payload_stateElements_3 = partialRound_inputBuffered_10_payload_stateElements_3;
  assign partialRound_bufferOut_3_payload_stateElements_4 = partialRound_inputBuffered_10_payload_stateElements_4;
  assign partialRound_bufferOut_3_payload_stateElements_5 = partialRound_inputBuffered_10_payload_stateElements_5;
  assign partialRound_bufferOut_3_payload_stateElements_6 = partialRound_inputBuffered_10_payload_stateElements_6;
  assign partialRound_bufferOut_3_payload_stateElements_7 = partialRound_inputBuffered_10_payload_stateElements_7;
  assign partialRound_bufferOut_3_payload_stateElements_8 = partialRound_inputBuffered_10_payload_stateElements_8;
  assign partialRound_bufferOut_3_payload_stateElements_9 = partialRound_inputBuffered_10_payload_stateElements_9;
  assign partialRound_bufferOut_3_payload_stateElements_10 = partialRound_inputBuffered_10_payload_stateElements_10;
  assign partialRound_bufferOut_3_payload_stateElements_11 = partialRound_inputBuffered_10_payload_stateElements_11;
  assign _zz_partialRound_bufferOutMuxed_valid = (partialRound_bufferOut_1_valid || partialRound_bufferOut_3_valid);
  assign _zz_partialRound_bufferOutMuxed_valid_1 = (partialRound_bufferOut_2_valid || partialRound_bufferOut_3_valid);
  assign _zz_partialRound_bufferOutMuxed_valid_2 = {_zz_partialRound_bufferOutMuxed_valid_1,_zz_partialRound_bufferOutMuxed_valid};
  assign partialRound_bufferOutMuxed_valid = _zz_partialRound_bufferOutMuxed_valid_3;
  assign partialRound_bufferOutMuxed_payload_isFull = _zz_partialRound_bufferOutMuxed_payload_isFull;
  assign partialRound_bufferOutMuxed_payload_fullRound = _zz_partialRound_bufferOutMuxed_payload_fullRound;
  assign partialRound_bufferOutMuxed_payload_partialRound = _zz_partialRound_bufferOutMuxed_payload_partialRound;
  assign partialRound_bufferOutMuxed_payload_stateSize = _zz_partialRound_bufferOutMuxed_payload_stateSize;
  assign partialRound_bufferOutMuxed_payload_stateID = _zz_partialRound_bufferOutMuxed_payload_stateID;
  assign partialRound_bufferOutMuxed_payload_stateElements_0 = _zz_partialRound_bufferOutMuxed_payload_stateElements_0;
  assign partialRound_bufferOutMuxed_payload_stateElements_1 = _zz_partialRound_bufferOutMuxed_payload_stateElements_1;
  assign partialRound_bufferOutMuxed_payload_stateElements_2 = _zz_partialRound_bufferOutMuxed_payload_stateElements_2;
  assign partialRound_bufferOutMuxed_payload_stateElements_3 = _zz_partialRound_bufferOutMuxed_payload_stateElements_3;
  assign partialRound_bufferOutMuxed_payload_stateElements_4 = _zz_partialRound_bufferOutMuxed_payload_stateElements_4;
  assign partialRound_bufferOutMuxed_payload_stateElements_5 = _zz_partialRound_bufferOutMuxed_payload_stateElements_5;
  assign partialRound_bufferOutMuxed_payload_stateElements_6 = _zz_partialRound_bufferOutMuxed_payload_stateElements_6;
  assign partialRound_bufferOutMuxed_payload_stateElements_7 = _zz_partialRound_bufferOutMuxed_payload_stateElements_7;
  assign partialRound_bufferOutMuxed_payload_stateElements_8 = _zz_partialRound_bufferOutMuxed_payload_stateElements_8;
  assign partialRound_bufferOutMuxed_payload_stateElements_9 = _zz_partialRound_bufferOutMuxed_payload_stateElements_9;
  assign partialRound_bufferOutMuxed_payload_stateElements_10 = _zz_partialRound_bufferOutMuxed_payload_stateElements_10;
  assign partialRound_bufferOutMuxed_payload_stateElements_11 = _zz_partialRound_bufferOutMuxed_payload_stateElements_11;
  assign when_MDSMatrixAdders_l67 = (partialRound_bufferOutMuxed_valid && (4'b0101 < partialRound_bufferOutMuxed_payload_stateSize));
  assign partialRound_bufferOutMuxed_takeWhen_valid = (partialRound_bufferOutMuxed_valid && (! partialRound_partialFlag));
  assign partialRound_bufferOutMuxed_takeWhen_payload_isFull = partialRound_bufferOutMuxed_payload_isFull;
  assign partialRound_bufferOutMuxed_takeWhen_payload_fullRound = partialRound_bufferOutMuxed_payload_fullRound;
  assign partialRound_bufferOutMuxed_takeWhen_payload_partialRound = partialRound_bufferOutMuxed_payload_partialRound;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateSize = partialRound_bufferOutMuxed_payload_stateSize;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateID = partialRound_bufferOutMuxed_payload_stateID;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_0 = partialRound_bufferOutMuxed_payload_stateElements_0;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_1 = partialRound_bufferOutMuxed_payload_stateElements_1;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_2 = partialRound_bufferOutMuxed_payload_stateElements_2;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_3 = partialRound_bufferOutMuxed_payload_stateElements_3;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_4 = partialRound_bufferOutMuxed_payload_stateElements_4;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_5 = partialRound_bufferOutMuxed_payload_stateElements_5;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_6 = partialRound_bufferOutMuxed_payload_stateElements_6;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_7 = partialRound_bufferOutMuxed_payload_stateElements_7;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_8 = partialRound_bufferOutMuxed_payload_stateElements_8;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_9 = partialRound_bufferOutMuxed_payload_stateElements_9;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_10 = partialRound_bufferOutMuxed_payload_stateElements_10;
  assign partialRound_bufferOutMuxed_takeWhen_payload_stateElements_11 = partialRound_bufferOutMuxed_payload_stateElements_11;
  always @(*) begin
    _zz_partialRound_adderTreeInput_payload_1 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_1 : partialRound_tempInput_payload_stateElements_1);
    if(when_MDSMatrixAdders_l75) begin
      _zz_partialRound_adderTreeInput_payload_1 = 255'h0;
    end else begin
      if(when_MDSMatrixAdders_l77) begin
        _zz_partialRound_adderTreeInput_payload_1 = 255'h0;
      end
    end
  end

  always @(*) begin
    _zz_partialRound_adderTreeInput_payload_2 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_2 : partialRound_tempInput_payload_stateElements_2);
    if(when_MDSMatrixAdders_l75) begin
      _zz_partialRound_adderTreeInput_payload_2 = 255'h0;
    end else begin
      if(when_MDSMatrixAdders_l77) begin
        _zz_partialRound_adderTreeInput_payload_2 = 255'h0;
      end
    end
  end

  always @(*) begin
    _zz_partialRound_adderTreeInput_payload_3 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_3 : partialRound_tempInput_payload_stateElements_3);
    if(!when_MDSMatrixAdders_l75) begin
      if(when_MDSMatrixAdders_l77) begin
        _zz_partialRound_adderTreeInput_payload_3 = 255'h0;
      end
    end
  end

  always @(*) begin
    _zz_partialRound_adderTreeInput_payload_4 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_4 : partialRound_tempInput_payload_stateElements_4);
    if(!when_MDSMatrixAdders_l75) begin
      if(when_MDSMatrixAdders_l77) begin
        _zz_partialRound_adderTreeInput_payload_4 = 255'h0;
      end
    end
  end

  assign when_MDSMatrixAdders_l75 = (partialRound_tempInput_payload_stateSize == 4'b0011);
  assign when_MDSMatrixAdders_l77 = (partialRound_tempInput_payload_stateSize == 4'b0101);
  assign partialRound_adderTreeInput_valid = partialRound_tempInput_valid;
  assign partialRound_adderTreeInput_payload_0 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_0 : partialRound_tempInput_payload_stateElements_0);
  assign partialRound_adderTreeInput_payload_1 = _zz_partialRound_adderTreeInput_payload_1;
  assign partialRound_adderTreeInput_payload_2 = _zz_partialRound_adderTreeInput_payload_2;
  assign partialRound_adderTreeInput_payload_3 = _zz_partialRound_adderTreeInput_payload_3;
  assign partialRound_adderTreeInput_payload_4 = _zz_partialRound_adderTreeInput_payload_4;
  assign partialRound_adderTreeInput_payload_5 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_5 : partialRound_tempInput_payload_stateElements_5);
  assign partialRound_adderTreeInput_payload_6 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_6 : partialRound_tempInput_payload_stateElements_6);
  assign partialRound_adderTreeInput_payload_7 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_7 : partialRound_tempInput_payload_stateElements_7);
  assign partialRound_adderTreeInput_payload_8 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_8 : partialRound_tempInput_payload_stateElements_8);
  assign partialRound_adderTreeInput_payload_9 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_9 : partialRound_tempInput_payload_stateElements_9);
  assign partialRound_adderTreeInput_payload_10 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_10 : partialRound_tempInput_payload_stateElements_10);
  assign partialRound_adderTreeInput_payload_11 = (partialRound_partialFlag ? partialRound_bufferOutMuxed_payload_stateElements_11 : partialRound_tempInput_payload_stateElements_11);
  always @(*) begin
    _zz_partialRound_output_payload_stateElements_0 = partialRound_contextDelayed_payload_stateElements_0;
    _zz_partialRound_output_payload_stateElements_0 = adderTree_1_io_output_payload;
  end

  always @(*) begin
    _zz_partialRound_output_payload_stateElements_3 = partialRound_contextDelayed_payload_stateElements_3;
    if(when_MDSMatrixAdders_l91) begin
      _zz_partialRound_output_payload_stateElements_3 = 255'h0;
    end
  end

  always @(*) begin
    _zz_partialRound_output_payload_stateElements_4 = partialRound_contextDelayed_payload_stateElements_4;
    if(when_MDSMatrixAdders_l91) begin
      _zz_partialRound_output_payload_stateElements_4 = 255'h0;
    end
  end

  always @(*) begin
    _zz_partialRound_output_payload_stateElements_5 = partialRound_contextDelayed_payload_stateElements_5;
    if(when_MDSMatrixAdders_l94) begin
      _zz_partialRound_output_payload_stateElements_5 = 255'h0;
    end
  end

  always @(*) begin
    _zz_partialRound_output_payload_stateElements_6 = partialRound_contextDelayed_payload_stateElements_6;
    if(when_MDSMatrixAdders_l94) begin
      _zz_partialRound_output_payload_stateElements_6 = 255'h0;
    end
  end

  always @(*) begin
    _zz_partialRound_output_payload_stateElements_7 = partialRound_contextDelayed_payload_stateElements_7;
    if(when_MDSMatrixAdders_l94) begin
      _zz_partialRound_output_payload_stateElements_7 = 255'h0;
    end
  end

  always @(*) begin
    _zz_partialRound_output_payload_stateElements_8 = partialRound_contextDelayed_payload_stateElements_8;
    if(when_MDSMatrixAdders_l94) begin
      _zz_partialRound_output_payload_stateElements_8 = 255'h0;
    end
  end

  assign when_MDSMatrixAdders_l91 = (partialRound_contextDelayed_payload_stateSize == 4'b0011);
  assign when_MDSMatrixAdders_l94 = (partialRound_contextDelayed_payload_stateSize == 4'b0101);
  assign fullRound_input_valid = (io_input_valid && io_input_payload_isFull);
  assign fullRound_input_payload_isFull = io_input_payload_isFull;
  assign fullRound_input_payload_fullRound = io_input_payload_fullRound;
  assign fullRound_input_payload_partialRound = io_input_payload_partialRound;
  assign fullRound_input_payload_stateSize = io_input_payload_stateSize;
  assign fullRound_input_payload_stateID = io_input_payload_stateID;
  assign fullRound_input_payload_stateElements_0 = io_input_payload_stateElements_0;
  assign fullRound_input_payload_stateElements_1 = io_input_payload_stateElements_1;
  assign fullRound_input_payload_stateElements_2 = io_input_payload_stateElements_2;
  assign fullRound_input_payload_stateElements_3 = io_input_payload_stateElements_3;
  assign fullRound_input_payload_stateElements_4 = io_input_payload_stateElements_4;
  assign fullRound_input_payload_stateElements_5 = io_input_payload_stateElements_5;
  assign fullRound_input_payload_stateElements_6 = io_input_payload_stateElements_6;
  assign fullRound_input_payload_stateElements_7 = io_input_payload_stateElements_7;
  assign fullRound_input_payload_stateElements_8 = io_input_payload_stateElements_8;
  assign fullRound_input_payload_stateElements_9 = io_input_payload_stateElements_9;
  assign fullRound_input_payload_stateElements_10 = io_input_payload_stateElements_10;
  assign fullRound_input_payload_stateElements_11 = io_input_payload_stateElements_11;
  assign fullRound_adderTreeInput_valid = fullRound_shiftMat_io_output_valid;
  assign fullRound_adderTreeInput_payload_0 = fullRound_shiftMat_io_output_payload_stateElements_0;
  assign fullRound_adderTreeInput_payload_1 = fullRound_shiftMat_io_output_payload_stateElements_1;
  assign fullRound_adderTreeInput_payload_2 = fullRound_shiftMat_io_output_payload_stateElements_2;
  assign fullRound_adderTreeInput_payload_3 = fullRound_shiftMat_io_output_payload_stateElements_3;
  assign fullRound_adderTreeInput_payload_4 = fullRound_shiftMat_io_output_payload_stateElements_4;
  assign fullRound_adderTreeInput_payload_5 = fullRound_shiftMat_io_output_payload_stateElements_5;
  assign fullRound_adderTreeInput_payload_6 = fullRound_shiftMat_io_output_payload_stateElements_6;
  assign fullRound_adderTreeInput_payload_7 = fullRound_shiftMat_io_output_payload_stateElements_7;
  assign fullRound_adderTreeInput_payload_8 = fullRound_shiftMat_io_output_payload_stateElements_8;
  assign fullRound_adderTreeInput_payload_9 = fullRound_shiftMat_io_output_payload_stateElements_9;
  assign fullRound_adderTreeInput_payload_10 = fullRound_shiftMat_io_output_payload_stateElements_10;
  assign fullRound_adderTreeInput_payload_11 = fullRound_shiftMat_io_output_payload_stateElements_11;
  assign fullRound_addContext_valid = fullRound_shiftMat_io_output_valid;
  assign fullRound_addContext_payload_isFull = fullRound_shiftMat_io_output_payload_isFull;
  assign fullRound_addContext_payload_fullRound = fullRound_shiftMat_io_output_payload_fullRound;
  assign fullRound_addContext_payload_partialRound = fullRound_shiftMat_io_output_payload_partialRound;
  assign fullRound_addContext_payload_stateSize = fullRound_shiftMat_io_output_payload_stateSize;
  assign fullRound_addContext_payload_stateID = fullRound_shiftMat_io_output_payload_stateID;
  assign fullRound_deserialization_wantExit = 1'b0;
  always @(*) begin
    fullRound_deserialization_wantStart = 1'b0;
    case(fullRound_deserialization_stateReg)
      fullRound_deserialization_enumDef_IDLE : begin
      end
      fullRound_deserialization_enumDef_BUSY : begin
      end
      fullRound_deserialization_enumDef_DONE : begin
      end
      default : begin
        fullRound_deserialization_wantStart = 1'b1;
      end
    endcase
  end

  assign fullRound_deserialization_wantKill = 1'b0;
  assign fullRound_output_payload_isFull = fullRound_deserialization_tempOutput_isFull;
  assign fullRound_output_payload_fullRound = fullRound_deserialization_tempOutput_fullRound;
  assign fullRound_output_payload_partialRound = fullRound_deserialization_tempOutput_partialRound;
  assign fullRound_output_payload_stateSize = fullRound_deserialization_tempOutput_stateSize;
  assign fullRound_output_payload_stateID = fullRound_deserialization_tempOutput_stateID;
  assign fullRound_output_payload_stateElements_0 = fullRound_deserialization_tempOutput_stateElements_0;
  assign fullRound_output_payload_stateElements_1 = fullRound_deserialization_tempOutput_stateElements_1;
  assign fullRound_output_payload_stateElements_2 = fullRound_deserialization_tempOutput_stateElements_2;
  assign fullRound_output_payload_stateElements_3 = fullRound_deserialization_tempOutput_stateElements_3;
  assign fullRound_output_payload_stateElements_4 = fullRound_deserialization_tempOutput_stateElements_4;
  assign fullRound_output_payload_stateElements_5 = fullRound_deserialization_tempOutput_stateElements_5;
  assign fullRound_output_payload_stateElements_6 = fullRound_deserialization_tempOutput_stateElements_6;
  assign fullRound_output_payload_stateElements_7 = fullRound_deserialization_tempOutput_stateElements_7;
  assign fullRound_output_payload_stateElements_8 = fullRound_deserialization_tempOutput_stateElements_8;
  assign fullRound_output_payload_stateElements_9 = fullRound_deserialization_tempOutput_stateElements_9;
  assign fullRound_output_payload_stateElements_10 = fullRound_deserialization_tempOutput_stateElements_10;
  assign fullRound_output_payload_stateElements_11 = fullRound_deserialization_tempOutput_stateElements_11;
  always @(*) begin
    fullRound_output_valid = 1'b0;
    case(fullRound_deserialization_stateReg)
      fullRound_deserialization_enumDef_IDLE : begin
      end
      fullRound_deserialization_enumDef_BUSY : begin
      end
      fullRound_deserialization_enumDef_DONE : begin
        fullRound_output_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign fullRound_deserialization_adderTreeValid = (adderTree_1_io_output_valid && fullRound_addContextDelayed_valid);
  always @(*) begin
    adderTree_1_io_input_valid = fullRound_adderTreeInput_valid;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_valid = partialRound_adderTreeInput_valid;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_0 = fullRound_adderTreeInput_payload_0;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_0 = partialRound_adderTreeInput_payload_0;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_1 = fullRound_adderTreeInput_payload_1;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_1 = partialRound_adderTreeInput_payload_1;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_2 = fullRound_adderTreeInput_payload_2;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_2 = partialRound_adderTreeInput_payload_2;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_3 = fullRound_adderTreeInput_payload_3;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_3 = partialRound_adderTreeInput_payload_3;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_4 = fullRound_adderTreeInput_payload_4;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_4 = partialRound_adderTreeInput_payload_4;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_5 = fullRound_adderTreeInput_payload_5;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_5 = partialRound_adderTreeInput_payload_5;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_6 = fullRound_adderTreeInput_payload_6;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_6 = partialRound_adderTreeInput_payload_6;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_7 = fullRound_adderTreeInput_payload_7;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_7 = partialRound_adderTreeInput_payload_7;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_8 = fullRound_adderTreeInput_payload_8;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_8 = partialRound_adderTreeInput_payload_8;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_9 = fullRound_adderTreeInput_payload_9;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_9 = partialRound_adderTreeInput_payload_9;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_10 = fullRound_adderTreeInput_payload_10;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_10 = partialRound_adderTreeInput_payload_10;
    end
  end

  always @(*) begin
    adderTree_1_io_input_payload_11 = fullRound_adderTreeInput_payload_11;
    if(partialRound_adderTreeInput_valid) begin
      adderTree_1_io_input_payload_11 = partialRound_adderTreeInput_payload_11;
    end
  end

  always @(*) begin
    io_output_valid = fullRound_output_valid;
    if(partialRound_output_valid) begin
      io_output_valid = partialRound_output_valid;
    end
  end

  always @(*) begin
    io_output_payload_isFull = fullRound_output_payload_isFull;
    if(partialRound_output_valid) begin
      io_output_payload_isFull = partialRound_output_payload_isFull;
    end
  end

  always @(*) begin
    io_output_payload_fullRound = fullRound_output_payload_fullRound;
    if(partialRound_output_valid) begin
      io_output_payload_fullRound = partialRound_output_payload_fullRound;
    end
  end

  always @(*) begin
    io_output_payload_partialRound = fullRound_output_payload_partialRound;
    if(partialRound_output_valid) begin
      io_output_payload_partialRound = partialRound_output_payload_partialRound;
    end
  end

  always @(*) begin
    io_output_payload_stateSize = fullRound_output_payload_stateSize;
    if(partialRound_output_valid) begin
      io_output_payload_stateSize = partialRound_output_payload_stateSize;
    end
  end

  always @(*) begin
    io_output_payload_stateID = fullRound_output_payload_stateID;
    if(partialRound_output_valid) begin
      io_output_payload_stateID = partialRound_output_payload_stateID;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_0 = fullRound_output_payload_stateElements_0;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_0 = partialRound_output_payload_stateElements_0;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_1 = fullRound_output_payload_stateElements_1;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_1 = partialRound_output_payload_stateElements_1;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_2 = fullRound_output_payload_stateElements_2;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_2 = partialRound_output_payload_stateElements_2;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_3 = fullRound_output_payload_stateElements_3;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_3 = partialRound_output_payload_stateElements_3;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_4 = fullRound_output_payload_stateElements_4;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_4 = partialRound_output_payload_stateElements_4;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_5 = fullRound_output_payload_stateElements_5;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_5 = partialRound_output_payload_stateElements_5;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_6 = fullRound_output_payload_stateElements_6;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_6 = partialRound_output_payload_stateElements_6;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_7 = fullRound_output_payload_stateElements_7;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_7 = partialRound_output_payload_stateElements_7;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_8 = fullRound_output_payload_stateElements_8;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_8 = partialRound_output_payload_stateElements_8;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_9 = fullRound_output_payload_stateElements_9;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_9 = partialRound_output_payload_stateElements_9;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_10 = fullRound_output_payload_stateElements_10;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_10 = partialRound_output_payload_stateElements_10;
    end
  end

  always @(*) begin
    io_output_payload_stateElements_11 = fullRound_output_payload_stateElements_11;
    if(partialRound_output_valid) begin
      io_output_payload_stateElements_11 = partialRound_output_payload_stateElements_11;
    end
  end

  always @(*) begin
    fullRound_deserialization_stateNext = fullRound_deserialization_stateReg;
    case(fullRound_deserialization_stateReg)
      fullRound_deserialization_enumDef_IDLE : begin
        if(fullRound_deserialization_adderTreeValid) begin
          fullRound_deserialization_stateNext = fullRound_deserialization_enumDef_BUSY;
        end
      end
      fullRound_deserialization_enumDef_BUSY : begin
        if(fullRound_deserialization_adderTreeValid) begin
          if(when_MDSMatrixAdders_l147) begin
            fullRound_deserialization_stateNext = fullRound_deserialization_enumDef_DONE;
          end
        end
      end
      fullRound_deserialization_enumDef_DONE : begin
        if(fullRound_deserialization_adderTreeValid) begin
          fullRound_deserialization_stateNext = fullRound_deserialization_enumDef_BUSY;
        end else begin
          fullRound_deserialization_stateNext = fullRound_deserialization_enumDef_IDLE;
        end
      end
      default : begin
      end
    endcase
    if(fullRound_deserialization_wantStart) begin
      fullRound_deserialization_stateNext = fullRound_deserialization_enumDef_IDLE;
    end
    if(fullRound_deserialization_wantKill) begin
      fullRound_deserialization_stateNext = fullRound_deserialization_enumDef_BOOT;
    end
  end

  assign _zz_1 = ({15'd0,1'b1} <<< fullRound_deserialization_counter);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = _zz_1[3];
  assign _zz_6 = _zz_1[4];
  assign _zz_7 = _zz_1[5];
  assign _zz_8 = _zz_1[6];
  assign _zz_9 = _zz_1[7];
  assign _zz_10 = _zz_1[8];
  assign _zz_11 = _zz_1[9];
  assign _zz_12 = _zz_1[10];
  assign _zz_13 = _zz_1[11];
  assign when_MDSMatrixAdders_l147 = (_zz_when_MDSMatrixAdders_l147 == fullRound_deserialization_tempOutput_stateSize);
  assign when_StateMachine_l222 = ((fullRound_deserialization_stateReg == fullRound_deserialization_enumDef_BUSY) && (! (fullRound_deserialization_stateNext == fullRound_deserialization_enumDef_BUSY)));
  always @(posedge clk) begin
    if(!resetn) begin
      partialRound_input_regNext_valid <= 1'b0;
      partialRound_inputBuffered_0_regNext_valid <= 1'b0;
      partialRound_inputBuffered_1_regNext_valid <= 1'b0;
      partialRound_inputBuffered_2_regNext_valid <= 1'b0;
      partialRound_inputBuffered_3_regNext_valid <= 1'b0;
      partialRound_inputBuffered_4_regNext_valid <= 1'b0;
      partialRound_inputBuffered_5_regNext_valid <= 1'b0;
      partialRound_inputBuffered_6_regNext_valid <= 1'b0;
      partialRound_inputBuffered_7_regNext_valid <= 1'b0;
      partialRound_inputBuffered_8_regNext_valid <= 1'b0;
      partialRound_inputBuffered_9_regNext_valid <= 1'b0;
      partialRound_partialFlag <= 1'b0;
      partialRound_tempInput_valid <= 1'b0;
      partialRound_output_valid <= 1'b0;
      fullRound_deserialization_counter <= 4'b0000;
      fullRound_deserialization_tempOutput_stateElements_0 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_1 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_2 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_3 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_4 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_5 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_6 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_7 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_8 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_9 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_10 <= 255'h0;
      fullRound_deserialization_tempOutput_stateElements_11 <= 255'h0;
      fullRound_deserialization_stateReg <= fullRound_deserialization_enumDef_BOOT;
    end else begin
      partialRound_input_regNext_valid <= partialRound_input_valid;
      partialRound_inputBuffered_0_regNext_valid <= partialRound_inputBuffered_0_valid;
      partialRound_inputBuffered_1_regNext_valid <= partialRound_inputBuffered_1_valid;
      partialRound_inputBuffered_2_regNext_valid <= partialRound_inputBuffered_2_valid;
      partialRound_inputBuffered_3_regNext_valid <= partialRound_inputBuffered_3_valid;
      partialRound_inputBuffered_4_regNext_valid <= partialRound_inputBuffered_4_valid;
      partialRound_inputBuffered_5_regNext_valid <= partialRound_inputBuffered_5_valid;
      partialRound_inputBuffered_6_regNext_valid <= partialRound_inputBuffered_6_valid;
      partialRound_inputBuffered_7_regNext_valid <= partialRound_inputBuffered_7_valid;
      partialRound_inputBuffered_8_regNext_valid <= partialRound_inputBuffered_8_valid;
      partialRound_inputBuffered_9_regNext_valid <= partialRound_inputBuffered_9_valid;
      if(when_MDSMatrixAdders_l67) begin
        partialRound_partialFlag <= (! partialRound_partialFlag);
      end
      partialRound_tempInput_valid <= partialRound_bufferOutMuxed_takeWhen_valid;
      partialRound_output_valid <= (adderTree_1_io_output_valid && partialRound_contextDelayed_valid);
      fullRound_deserialization_stateReg <= fullRound_deserialization_stateNext;
      case(fullRound_deserialization_stateReg)
        fullRound_deserialization_enumDef_IDLE : begin
          if(fullRound_deserialization_adderTreeValid) begin
            if(_zz_2) begin
              fullRound_deserialization_tempOutput_stateElements_0 <= adderTree_1_io_output_payload;
            end
            if(_zz_3) begin
              fullRound_deserialization_tempOutput_stateElements_1 <= adderTree_1_io_output_payload;
            end
            if(_zz_4) begin
              fullRound_deserialization_tempOutput_stateElements_2 <= adderTree_1_io_output_payload;
            end
            if(_zz_5) begin
              fullRound_deserialization_tempOutput_stateElements_3 <= adderTree_1_io_output_payload;
            end
            if(_zz_6) begin
              fullRound_deserialization_tempOutput_stateElements_4 <= adderTree_1_io_output_payload;
            end
            if(_zz_7) begin
              fullRound_deserialization_tempOutput_stateElements_5 <= adderTree_1_io_output_payload;
            end
            if(_zz_8) begin
              fullRound_deserialization_tempOutput_stateElements_6 <= adderTree_1_io_output_payload;
            end
            if(_zz_9) begin
              fullRound_deserialization_tempOutput_stateElements_7 <= adderTree_1_io_output_payload;
            end
            if(_zz_10) begin
              fullRound_deserialization_tempOutput_stateElements_8 <= adderTree_1_io_output_payload;
            end
            if(_zz_11) begin
              fullRound_deserialization_tempOutput_stateElements_9 <= adderTree_1_io_output_payload;
            end
            if(_zz_12) begin
              fullRound_deserialization_tempOutput_stateElements_10 <= adderTree_1_io_output_payload;
            end
            if(_zz_13) begin
              fullRound_deserialization_tempOutput_stateElements_11 <= adderTree_1_io_output_payload;
            end
            fullRound_deserialization_counter <= (fullRound_deserialization_counter + 4'b0001);
          end
        end
        fullRound_deserialization_enumDef_BUSY : begin
          if(fullRound_deserialization_adderTreeValid) begin
            if(_zz_2) begin
              fullRound_deserialization_tempOutput_stateElements_0 <= adderTree_1_io_output_payload;
            end
            if(_zz_3) begin
              fullRound_deserialization_tempOutput_stateElements_1 <= adderTree_1_io_output_payload;
            end
            if(_zz_4) begin
              fullRound_deserialization_tempOutput_stateElements_2 <= adderTree_1_io_output_payload;
            end
            if(_zz_5) begin
              fullRound_deserialization_tempOutput_stateElements_3 <= adderTree_1_io_output_payload;
            end
            if(_zz_6) begin
              fullRound_deserialization_tempOutput_stateElements_4 <= adderTree_1_io_output_payload;
            end
            if(_zz_7) begin
              fullRound_deserialization_tempOutput_stateElements_5 <= adderTree_1_io_output_payload;
            end
            if(_zz_8) begin
              fullRound_deserialization_tempOutput_stateElements_6 <= adderTree_1_io_output_payload;
            end
            if(_zz_9) begin
              fullRound_deserialization_tempOutput_stateElements_7 <= adderTree_1_io_output_payload;
            end
            if(_zz_10) begin
              fullRound_deserialization_tempOutput_stateElements_8 <= adderTree_1_io_output_payload;
            end
            if(_zz_11) begin
              fullRound_deserialization_tempOutput_stateElements_9 <= adderTree_1_io_output_payload;
            end
            if(_zz_12) begin
              fullRound_deserialization_tempOutput_stateElements_10 <= adderTree_1_io_output_payload;
            end
            if(_zz_13) begin
              fullRound_deserialization_tempOutput_stateElements_11 <= adderTree_1_io_output_payload;
            end
            if(!when_MDSMatrixAdders_l147) begin
              fullRound_deserialization_counter <= (fullRound_deserialization_counter + 4'b0001);
            end
          end
        end
        fullRound_deserialization_enumDef_DONE : begin
          if(fullRound_deserialization_adderTreeValid) begin
            if(_zz_2) begin
              fullRound_deserialization_tempOutput_stateElements_0 <= adderTree_1_io_output_payload;
            end
            if(_zz_3) begin
              fullRound_deserialization_tempOutput_stateElements_1 <= adderTree_1_io_output_payload;
            end
            if(_zz_4) begin
              fullRound_deserialization_tempOutput_stateElements_2 <= adderTree_1_io_output_payload;
            end
            if(_zz_5) begin
              fullRound_deserialization_tempOutput_stateElements_3 <= adderTree_1_io_output_payload;
            end
            if(_zz_6) begin
              fullRound_deserialization_tempOutput_stateElements_4 <= adderTree_1_io_output_payload;
            end
            if(_zz_7) begin
              fullRound_deserialization_tempOutput_stateElements_5 <= adderTree_1_io_output_payload;
            end
            if(_zz_8) begin
              fullRound_deserialization_tempOutput_stateElements_6 <= adderTree_1_io_output_payload;
            end
            if(_zz_9) begin
              fullRound_deserialization_tempOutput_stateElements_7 <= adderTree_1_io_output_payload;
            end
            if(_zz_10) begin
              fullRound_deserialization_tempOutput_stateElements_8 <= adderTree_1_io_output_payload;
            end
            if(_zz_11) begin
              fullRound_deserialization_tempOutput_stateElements_9 <= adderTree_1_io_output_payload;
            end
            if(_zz_12) begin
              fullRound_deserialization_tempOutput_stateElements_10 <= adderTree_1_io_output_payload;
            end
            if(_zz_13) begin
              fullRound_deserialization_tempOutput_stateElements_11 <= adderTree_1_io_output_payload;
            end
            fullRound_deserialization_counter <= (fullRound_deserialization_counter + 4'b0001);
          end
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l222) begin
        fullRound_deserialization_counter <= 4'b0000;
      end
    end
  end

  always @(posedge clk) begin
    partialRound_input_regNext_payload_isFull <= partialRound_input_payload_isFull;
    partialRound_input_regNext_payload_fullRound <= partialRound_input_payload_fullRound;
    partialRound_input_regNext_payload_partialRound <= partialRound_input_payload_partialRound;
    partialRound_input_regNext_payload_stateSize <= partialRound_input_payload_stateSize;
    partialRound_input_regNext_payload_stateID <= partialRound_input_payload_stateID;
    partialRound_input_regNext_payload_stateElements_0 <= partialRound_input_payload_stateElements_0;
    partialRound_input_regNext_payload_stateElements_1 <= partialRound_input_payload_stateElements_1;
    partialRound_input_regNext_payload_stateElements_2 <= partialRound_input_payload_stateElements_2;
    partialRound_input_regNext_payload_stateElements_3 <= partialRound_input_payload_stateElements_3;
    partialRound_input_regNext_payload_stateElements_4 <= partialRound_input_payload_stateElements_4;
    partialRound_input_regNext_payload_stateElements_5 <= partialRound_input_payload_stateElements_5;
    partialRound_input_regNext_payload_stateElements_6 <= partialRound_input_payload_stateElements_6;
    partialRound_input_regNext_payload_stateElements_7 <= partialRound_input_payload_stateElements_7;
    partialRound_input_regNext_payload_stateElements_8 <= partialRound_input_payload_stateElements_8;
    partialRound_input_regNext_payload_stateElements_9 <= partialRound_input_payload_stateElements_9;
    partialRound_input_regNext_payload_stateElements_10 <= partialRound_input_payload_stateElements_10;
    partialRound_input_regNext_payload_stateElements_11 <= partialRound_input_payload_stateElements_11;
    partialRound_inputBuffered_0_regNext_payload_isFull <= partialRound_inputBuffered_0_payload_isFull;
    partialRound_inputBuffered_0_regNext_payload_fullRound <= partialRound_inputBuffered_0_payload_fullRound;
    partialRound_inputBuffered_0_regNext_payload_partialRound <= partialRound_inputBuffered_0_payload_partialRound;
    partialRound_inputBuffered_0_regNext_payload_stateSize <= partialRound_inputBuffered_0_payload_stateSize;
    partialRound_inputBuffered_0_regNext_payload_stateID <= partialRound_inputBuffered_0_payload_stateID;
    partialRound_inputBuffered_0_regNext_payload_stateElements_0 <= partialRound_inputBuffered_0_payload_stateElements_0;
    partialRound_inputBuffered_0_regNext_payload_stateElements_1 <= partialRound_inputBuffered_0_payload_stateElements_1;
    partialRound_inputBuffered_0_regNext_payload_stateElements_2 <= partialRound_inputBuffered_0_payload_stateElements_2;
    partialRound_inputBuffered_0_regNext_payload_stateElements_3 <= partialRound_inputBuffered_0_payload_stateElements_3;
    partialRound_inputBuffered_0_regNext_payload_stateElements_4 <= partialRound_inputBuffered_0_payload_stateElements_4;
    partialRound_inputBuffered_0_regNext_payload_stateElements_5 <= partialRound_inputBuffered_0_payload_stateElements_5;
    partialRound_inputBuffered_0_regNext_payload_stateElements_6 <= partialRound_inputBuffered_0_payload_stateElements_6;
    partialRound_inputBuffered_0_regNext_payload_stateElements_7 <= partialRound_inputBuffered_0_payload_stateElements_7;
    partialRound_inputBuffered_0_regNext_payload_stateElements_8 <= partialRound_inputBuffered_0_payload_stateElements_8;
    partialRound_inputBuffered_0_regNext_payload_stateElements_9 <= partialRound_inputBuffered_0_payload_stateElements_9;
    partialRound_inputBuffered_0_regNext_payload_stateElements_10 <= partialRound_inputBuffered_0_payload_stateElements_10;
    partialRound_inputBuffered_0_regNext_payload_stateElements_11 <= partialRound_inputBuffered_0_payload_stateElements_11;
    partialRound_inputBuffered_1_regNext_payload_isFull <= partialRound_inputBuffered_1_payload_isFull;
    partialRound_inputBuffered_1_regNext_payload_fullRound <= partialRound_inputBuffered_1_payload_fullRound;
    partialRound_inputBuffered_1_regNext_payload_partialRound <= partialRound_inputBuffered_1_payload_partialRound;
    partialRound_inputBuffered_1_regNext_payload_stateSize <= partialRound_inputBuffered_1_payload_stateSize;
    partialRound_inputBuffered_1_regNext_payload_stateID <= partialRound_inputBuffered_1_payload_stateID;
    partialRound_inputBuffered_1_regNext_payload_stateElements_0 <= partialRound_inputBuffered_1_payload_stateElements_0;
    partialRound_inputBuffered_1_regNext_payload_stateElements_1 <= partialRound_inputBuffered_1_payload_stateElements_1;
    partialRound_inputBuffered_1_regNext_payload_stateElements_2 <= partialRound_inputBuffered_1_payload_stateElements_2;
    partialRound_inputBuffered_1_regNext_payload_stateElements_3 <= partialRound_inputBuffered_1_payload_stateElements_3;
    partialRound_inputBuffered_1_regNext_payload_stateElements_4 <= partialRound_inputBuffered_1_payload_stateElements_4;
    partialRound_inputBuffered_1_regNext_payload_stateElements_5 <= partialRound_inputBuffered_1_payload_stateElements_5;
    partialRound_inputBuffered_1_regNext_payload_stateElements_6 <= partialRound_inputBuffered_1_payload_stateElements_6;
    partialRound_inputBuffered_1_regNext_payload_stateElements_7 <= partialRound_inputBuffered_1_payload_stateElements_7;
    partialRound_inputBuffered_1_regNext_payload_stateElements_8 <= partialRound_inputBuffered_1_payload_stateElements_8;
    partialRound_inputBuffered_1_regNext_payload_stateElements_9 <= partialRound_inputBuffered_1_payload_stateElements_9;
    partialRound_inputBuffered_1_regNext_payload_stateElements_10 <= partialRound_inputBuffered_1_payload_stateElements_10;
    partialRound_inputBuffered_1_regNext_payload_stateElements_11 <= partialRound_inputBuffered_1_payload_stateElements_11;
    partialRound_inputBuffered_2_regNext_payload_isFull <= partialRound_inputBuffered_2_payload_isFull;
    partialRound_inputBuffered_2_regNext_payload_fullRound <= partialRound_inputBuffered_2_payload_fullRound;
    partialRound_inputBuffered_2_regNext_payload_partialRound <= partialRound_inputBuffered_2_payload_partialRound;
    partialRound_inputBuffered_2_regNext_payload_stateSize <= partialRound_inputBuffered_2_payload_stateSize;
    partialRound_inputBuffered_2_regNext_payload_stateID <= partialRound_inputBuffered_2_payload_stateID;
    partialRound_inputBuffered_2_regNext_payload_stateElements_0 <= partialRound_inputBuffered_2_payload_stateElements_0;
    partialRound_inputBuffered_2_regNext_payload_stateElements_1 <= partialRound_inputBuffered_2_payload_stateElements_1;
    partialRound_inputBuffered_2_regNext_payload_stateElements_2 <= partialRound_inputBuffered_2_payload_stateElements_2;
    partialRound_inputBuffered_2_regNext_payload_stateElements_3 <= partialRound_inputBuffered_2_payload_stateElements_3;
    partialRound_inputBuffered_2_regNext_payload_stateElements_4 <= partialRound_inputBuffered_2_payload_stateElements_4;
    partialRound_inputBuffered_2_regNext_payload_stateElements_5 <= partialRound_inputBuffered_2_payload_stateElements_5;
    partialRound_inputBuffered_2_regNext_payload_stateElements_6 <= partialRound_inputBuffered_2_payload_stateElements_6;
    partialRound_inputBuffered_2_regNext_payload_stateElements_7 <= partialRound_inputBuffered_2_payload_stateElements_7;
    partialRound_inputBuffered_2_regNext_payload_stateElements_8 <= partialRound_inputBuffered_2_payload_stateElements_8;
    partialRound_inputBuffered_2_regNext_payload_stateElements_9 <= partialRound_inputBuffered_2_payload_stateElements_9;
    partialRound_inputBuffered_2_regNext_payload_stateElements_10 <= partialRound_inputBuffered_2_payload_stateElements_10;
    partialRound_inputBuffered_2_regNext_payload_stateElements_11 <= partialRound_inputBuffered_2_payload_stateElements_11;
    partialRound_inputBuffered_3_regNext_payload_isFull <= partialRound_inputBuffered_3_payload_isFull;
    partialRound_inputBuffered_3_regNext_payload_fullRound <= partialRound_inputBuffered_3_payload_fullRound;
    partialRound_inputBuffered_3_regNext_payload_partialRound <= partialRound_inputBuffered_3_payload_partialRound;
    partialRound_inputBuffered_3_regNext_payload_stateSize <= partialRound_inputBuffered_3_payload_stateSize;
    partialRound_inputBuffered_3_regNext_payload_stateID <= partialRound_inputBuffered_3_payload_stateID;
    partialRound_inputBuffered_3_regNext_payload_stateElements_0 <= partialRound_inputBuffered_3_payload_stateElements_0;
    partialRound_inputBuffered_3_regNext_payload_stateElements_1 <= partialRound_inputBuffered_3_payload_stateElements_1;
    partialRound_inputBuffered_3_regNext_payload_stateElements_2 <= partialRound_inputBuffered_3_payload_stateElements_2;
    partialRound_inputBuffered_3_regNext_payload_stateElements_3 <= partialRound_inputBuffered_3_payload_stateElements_3;
    partialRound_inputBuffered_3_regNext_payload_stateElements_4 <= partialRound_inputBuffered_3_payload_stateElements_4;
    partialRound_inputBuffered_3_regNext_payload_stateElements_5 <= partialRound_inputBuffered_3_payload_stateElements_5;
    partialRound_inputBuffered_3_regNext_payload_stateElements_6 <= partialRound_inputBuffered_3_payload_stateElements_6;
    partialRound_inputBuffered_3_regNext_payload_stateElements_7 <= partialRound_inputBuffered_3_payload_stateElements_7;
    partialRound_inputBuffered_3_regNext_payload_stateElements_8 <= partialRound_inputBuffered_3_payload_stateElements_8;
    partialRound_inputBuffered_3_regNext_payload_stateElements_9 <= partialRound_inputBuffered_3_payload_stateElements_9;
    partialRound_inputBuffered_3_regNext_payload_stateElements_10 <= partialRound_inputBuffered_3_payload_stateElements_10;
    partialRound_inputBuffered_3_regNext_payload_stateElements_11 <= partialRound_inputBuffered_3_payload_stateElements_11;
    partialRound_inputBuffered_4_regNext_payload_isFull <= partialRound_inputBuffered_4_payload_isFull;
    partialRound_inputBuffered_4_regNext_payload_fullRound <= partialRound_inputBuffered_4_payload_fullRound;
    partialRound_inputBuffered_4_regNext_payload_partialRound <= partialRound_inputBuffered_4_payload_partialRound;
    partialRound_inputBuffered_4_regNext_payload_stateSize <= partialRound_inputBuffered_4_payload_stateSize;
    partialRound_inputBuffered_4_regNext_payload_stateID <= partialRound_inputBuffered_4_payload_stateID;
    partialRound_inputBuffered_4_regNext_payload_stateElements_0 <= partialRound_inputBuffered_4_payload_stateElements_0;
    partialRound_inputBuffered_4_regNext_payload_stateElements_1 <= partialRound_inputBuffered_4_payload_stateElements_1;
    partialRound_inputBuffered_4_regNext_payload_stateElements_2 <= partialRound_inputBuffered_4_payload_stateElements_2;
    partialRound_inputBuffered_4_regNext_payload_stateElements_3 <= partialRound_inputBuffered_4_payload_stateElements_3;
    partialRound_inputBuffered_4_regNext_payload_stateElements_4 <= partialRound_inputBuffered_4_payload_stateElements_4;
    partialRound_inputBuffered_4_regNext_payload_stateElements_5 <= partialRound_inputBuffered_4_payload_stateElements_5;
    partialRound_inputBuffered_4_regNext_payload_stateElements_6 <= partialRound_inputBuffered_4_payload_stateElements_6;
    partialRound_inputBuffered_4_regNext_payload_stateElements_7 <= partialRound_inputBuffered_4_payload_stateElements_7;
    partialRound_inputBuffered_4_regNext_payload_stateElements_8 <= partialRound_inputBuffered_4_payload_stateElements_8;
    partialRound_inputBuffered_4_regNext_payload_stateElements_9 <= partialRound_inputBuffered_4_payload_stateElements_9;
    partialRound_inputBuffered_4_regNext_payload_stateElements_10 <= partialRound_inputBuffered_4_payload_stateElements_10;
    partialRound_inputBuffered_4_regNext_payload_stateElements_11 <= partialRound_inputBuffered_4_payload_stateElements_11;
    partialRound_inputBuffered_5_regNext_payload_isFull <= partialRound_inputBuffered_5_payload_isFull;
    partialRound_inputBuffered_5_regNext_payload_fullRound <= partialRound_inputBuffered_5_payload_fullRound;
    partialRound_inputBuffered_5_regNext_payload_partialRound <= partialRound_inputBuffered_5_payload_partialRound;
    partialRound_inputBuffered_5_regNext_payload_stateSize <= partialRound_inputBuffered_5_payload_stateSize;
    partialRound_inputBuffered_5_regNext_payload_stateID <= partialRound_inputBuffered_5_payload_stateID;
    partialRound_inputBuffered_5_regNext_payload_stateElements_0 <= partialRound_inputBuffered_5_payload_stateElements_0;
    partialRound_inputBuffered_5_regNext_payload_stateElements_1 <= partialRound_inputBuffered_5_payload_stateElements_1;
    partialRound_inputBuffered_5_regNext_payload_stateElements_2 <= partialRound_inputBuffered_5_payload_stateElements_2;
    partialRound_inputBuffered_5_regNext_payload_stateElements_3 <= partialRound_inputBuffered_5_payload_stateElements_3;
    partialRound_inputBuffered_5_regNext_payload_stateElements_4 <= partialRound_inputBuffered_5_payload_stateElements_4;
    partialRound_inputBuffered_5_regNext_payload_stateElements_5 <= partialRound_inputBuffered_5_payload_stateElements_5;
    partialRound_inputBuffered_5_regNext_payload_stateElements_6 <= partialRound_inputBuffered_5_payload_stateElements_6;
    partialRound_inputBuffered_5_regNext_payload_stateElements_7 <= partialRound_inputBuffered_5_payload_stateElements_7;
    partialRound_inputBuffered_5_regNext_payload_stateElements_8 <= partialRound_inputBuffered_5_payload_stateElements_8;
    partialRound_inputBuffered_5_regNext_payload_stateElements_9 <= partialRound_inputBuffered_5_payload_stateElements_9;
    partialRound_inputBuffered_5_regNext_payload_stateElements_10 <= partialRound_inputBuffered_5_payload_stateElements_10;
    partialRound_inputBuffered_5_regNext_payload_stateElements_11 <= partialRound_inputBuffered_5_payload_stateElements_11;
    partialRound_inputBuffered_6_regNext_payload_isFull <= partialRound_inputBuffered_6_payload_isFull;
    partialRound_inputBuffered_6_regNext_payload_fullRound <= partialRound_inputBuffered_6_payload_fullRound;
    partialRound_inputBuffered_6_regNext_payload_partialRound <= partialRound_inputBuffered_6_payload_partialRound;
    partialRound_inputBuffered_6_regNext_payload_stateSize <= partialRound_inputBuffered_6_payload_stateSize;
    partialRound_inputBuffered_6_regNext_payload_stateID <= partialRound_inputBuffered_6_payload_stateID;
    partialRound_inputBuffered_6_regNext_payload_stateElements_0 <= partialRound_inputBuffered_6_payload_stateElements_0;
    partialRound_inputBuffered_6_regNext_payload_stateElements_1 <= partialRound_inputBuffered_6_payload_stateElements_1;
    partialRound_inputBuffered_6_regNext_payload_stateElements_2 <= partialRound_inputBuffered_6_payload_stateElements_2;
    partialRound_inputBuffered_6_regNext_payload_stateElements_3 <= partialRound_inputBuffered_6_payload_stateElements_3;
    partialRound_inputBuffered_6_regNext_payload_stateElements_4 <= partialRound_inputBuffered_6_payload_stateElements_4;
    partialRound_inputBuffered_6_regNext_payload_stateElements_5 <= partialRound_inputBuffered_6_payload_stateElements_5;
    partialRound_inputBuffered_6_regNext_payload_stateElements_6 <= partialRound_inputBuffered_6_payload_stateElements_6;
    partialRound_inputBuffered_6_regNext_payload_stateElements_7 <= partialRound_inputBuffered_6_payload_stateElements_7;
    partialRound_inputBuffered_6_regNext_payload_stateElements_8 <= partialRound_inputBuffered_6_payload_stateElements_8;
    partialRound_inputBuffered_6_regNext_payload_stateElements_9 <= partialRound_inputBuffered_6_payload_stateElements_9;
    partialRound_inputBuffered_6_regNext_payload_stateElements_10 <= partialRound_inputBuffered_6_payload_stateElements_10;
    partialRound_inputBuffered_6_regNext_payload_stateElements_11 <= partialRound_inputBuffered_6_payload_stateElements_11;
    partialRound_inputBuffered_7_regNext_payload_isFull <= partialRound_inputBuffered_7_payload_isFull;
    partialRound_inputBuffered_7_regNext_payload_fullRound <= partialRound_inputBuffered_7_payload_fullRound;
    partialRound_inputBuffered_7_regNext_payload_partialRound <= partialRound_inputBuffered_7_payload_partialRound;
    partialRound_inputBuffered_7_regNext_payload_stateSize <= partialRound_inputBuffered_7_payload_stateSize;
    partialRound_inputBuffered_7_regNext_payload_stateID <= partialRound_inputBuffered_7_payload_stateID;
    partialRound_inputBuffered_7_regNext_payload_stateElements_0 <= partialRound_inputBuffered_7_payload_stateElements_0;
    partialRound_inputBuffered_7_regNext_payload_stateElements_1 <= partialRound_inputBuffered_7_payload_stateElements_1;
    partialRound_inputBuffered_7_regNext_payload_stateElements_2 <= partialRound_inputBuffered_7_payload_stateElements_2;
    partialRound_inputBuffered_7_regNext_payload_stateElements_3 <= partialRound_inputBuffered_7_payload_stateElements_3;
    partialRound_inputBuffered_7_regNext_payload_stateElements_4 <= partialRound_inputBuffered_7_payload_stateElements_4;
    partialRound_inputBuffered_7_regNext_payload_stateElements_5 <= partialRound_inputBuffered_7_payload_stateElements_5;
    partialRound_inputBuffered_7_regNext_payload_stateElements_6 <= partialRound_inputBuffered_7_payload_stateElements_6;
    partialRound_inputBuffered_7_regNext_payload_stateElements_7 <= partialRound_inputBuffered_7_payload_stateElements_7;
    partialRound_inputBuffered_7_regNext_payload_stateElements_8 <= partialRound_inputBuffered_7_payload_stateElements_8;
    partialRound_inputBuffered_7_regNext_payload_stateElements_9 <= partialRound_inputBuffered_7_payload_stateElements_9;
    partialRound_inputBuffered_7_regNext_payload_stateElements_10 <= partialRound_inputBuffered_7_payload_stateElements_10;
    partialRound_inputBuffered_7_regNext_payload_stateElements_11 <= partialRound_inputBuffered_7_payload_stateElements_11;
    partialRound_inputBuffered_8_regNext_payload_isFull <= partialRound_inputBuffered_8_payload_isFull;
    partialRound_inputBuffered_8_regNext_payload_fullRound <= partialRound_inputBuffered_8_payload_fullRound;
    partialRound_inputBuffered_8_regNext_payload_partialRound <= partialRound_inputBuffered_8_payload_partialRound;
    partialRound_inputBuffered_8_regNext_payload_stateSize <= partialRound_inputBuffered_8_payload_stateSize;
    partialRound_inputBuffered_8_regNext_payload_stateID <= partialRound_inputBuffered_8_payload_stateID;
    partialRound_inputBuffered_8_regNext_payload_stateElements_0 <= partialRound_inputBuffered_8_payload_stateElements_0;
    partialRound_inputBuffered_8_regNext_payload_stateElements_1 <= partialRound_inputBuffered_8_payload_stateElements_1;
    partialRound_inputBuffered_8_regNext_payload_stateElements_2 <= partialRound_inputBuffered_8_payload_stateElements_2;
    partialRound_inputBuffered_8_regNext_payload_stateElements_3 <= partialRound_inputBuffered_8_payload_stateElements_3;
    partialRound_inputBuffered_8_regNext_payload_stateElements_4 <= partialRound_inputBuffered_8_payload_stateElements_4;
    partialRound_inputBuffered_8_regNext_payload_stateElements_5 <= partialRound_inputBuffered_8_payload_stateElements_5;
    partialRound_inputBuffered_8_regNext_payload_stateElements_6 <= partialRound_inputBuffered_8_payload_stateElements_6;
    partialRound_inputBuffered_8_regNext_payload_stateElements_7 <= partialRound_inputBuffered_8_payload_stateElements_7;
    partialRound_inputBuffered_8_regNext_payload_stateElements_8 <= partialRound_inputBuffered_8_payload_stateElements_8;
    partialRound_inputBuffered_8_regNext_payload_stateElements_9 <= partialRound_inputBuffered_8_payload_stateElements_9;
    partialRound_inputBuffered_8_regNext_payload_stateElements_10 <= partialRound_inputBuffered_8_payload_stateElements_10;
    partialRound_inputBuffered_8_regNext_payload_stateElements_11 <= partialRound_inputBuffered_8_payload_stateElements_11;
    partialRound_inputBuffered_9_regNext_payload_isFull <= partialRound_inputBuffered_9_payload_isFull;
    partialRound_inputBuffered_9_regNext_payload_fullRound <= partialRound_inputBuffered_9_payload_fullRound;
    partialRound_inputBuffered_9_regNext_payload_partialRound <= partialRound_inputBuffered_9_payload_partialRound;
    partialRound_inputBuffered_9_regNext_payload_stateSize <= partialRound_inputBuffered_9_payload_stateSize;
    partialRound_inputBuffered_9_regNext_payload_stateID <= partialRound_inputBuffered_9_payload_stateID;
    partialRound_inputBuffered_9_regNext_payload_stateElements_0 <= partialRound_inputBuffered_9_payload_stateElements_0;
    partialRound_inputBuffered_9_regNext_payload_stateElements_1 <= partialRound_inputBuffered_9_payload_stateElements_1;
    partialRound_inputBuffered_9_regNext_payload_stateElements_2 <= partialRound_inputBuffered_9_payload_stateElements_2;
    partialRound_inputBuffered_9_regNext_payload_stateElements_3 <= partialRound_inputBuffered_9_payload_stateElements_3;
    partialRound_inputBuffered_9_regNext_payload_stateElements_4 <= partialRound_inputBuffered_9_payload_stateElements_4;
    partialRound_inputBuffered_9_regNext_payload_stateElements_5 <= partialRound_inputBuffered_9_payload_stateElements_5;
    partialRound_inputBuffered_9_regNext_payload_stateElements_6 <= partialRound_inputBuffered_9_payload_stateElements_6;
    partialRound_inputBuffered_9_regNext_payload_stateElements_7 <= partialRound_inputBuffered_9_payload_stateElements_7;
    partialRound_inputBuffered_9_regNext_payload_stateElements_8 <= partialRound_inputBuffered_9_payload_stateElements_8;
    partialRound_inputBuffered_9_regNext_payload_stateElements_9 <= partialRound_inputBuffered_9_payload_stateElements_9;
    partialRound_inputBuffered_9_regNext_payload_stateElements_10 <= partialRound_inputBuffered_9_payload_stateElements_10;
    partialRound_inputBuffered_9_regNext_payload_stateElements_11 <= partialRound_inputBuffered_9_payload_stateElements_11;
    partialRound_tempInput_payload_isFull <= partialRound_bufferOutMuxed_takeWhen_payload_isFull;
    partialRound_tempInput_payload_fullRound <= partialRound_bufferOutMuxed_takeWhen_payload_fullRound;
    partialRound_tempInput_payload_partialRound <= partialRound_bufferOutMuxed_takeWhen_payload_partialRound;
    partialRound_tempInput_payload_stateSize <= partialRound_bufferOutMuxed_takeWhen_payload_stateSize;
    partialRound_tempInput_payload_stateID <= partialRound_bufferOutMuxed_takeWhen_payload_stateID;
    partialRound_tempInput_payload_stateElements_0 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_0;
    partialRound_tempInput_payload_stateElements_1 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_1;
    partialRound_tempInput_payload_stateElements_2 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_2;
    partialRound_tempInput_payload_stateElements_3 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_3;
    partialRound_tempInput_payload_stateElements_4 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_4;
    partialRound_tempInput_payload_stateElements_5 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_5;
    partialRound_tempInput_payload_stateElements_6 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_6;
    partialRound_tempInput_payload_stateElements_7 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_7;
    partialRound_tempInput_payload_stateElements_8 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_8;
    partialRound_tempInput_payload_stateElements_9 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_9;
    partialRound_tempInput_payload_stateElements_10 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_10;
    partialRound_tempInput_payload_stateElements_11 <= partialRound_bufferOutMuxed_takeWhen_payload_stateElements_11;
    partialRound_tempInput_delay_1_valid <= partialRound_tempInput_valid;
    partialRound_tempInput_delay_1_payload_isFull <= partialRound_tempInput_payload_isFull;
    partialRound_tempInput_delay_1_payload_fullRound <= partialRound_tempInput_payload_fullRound;
    partialRound_tempInput_delay_1_payload_partialRound <= partialRound_tempInput_payload_partialRound;
    partialRound_tempInput_delay_1_payload_stateSize <= partialRound_tempInput_payload_stateSize;
    partialRound_tempInput_delay_1_payload_stateID <= partialRound_tempInput_payload_stateID;
    partialRound_tempInput_delay_1_payload_stateElements_0 <= partialRound_tempInput_payload_stateElements_0;
    partialRound_tempInput_delay_1_payload_stateElements_1 <= partialRound_tempInput_payload_stateElements_1;
    partialRound_tempInput_delay_1_payload_stateElements_2 <= partialRound_tempInput_payload_stateElements_2;
    partialRound_tempInput_delay_1_payload_stateElements_3 <= partialRound_tempInput_payload_stateElements_3;
    partialRound_tempInput_delay_1_payload_stateElements_4 <= partialRound_tempInput_payload_stateElements_4;
    partialRound_tempInput_delay_1_payload_stateElements_5 <= partialRound_tempInput_payload_stateElements_5;
    partialRound_tempInput_delay_1_payload_stateElements_6 <= partialRound_tempInput_payload_stateElements_6;
    partialRound_tempInput_delay_1_payload_stateElements_7 <= partialRound_tempInput_payload_stateElements_7;
    partialRound_tempInput_delay_1_payload_stateElements_8 <= partialRound_tempInput_payload_stateElements_8;
    partialRound_tempInput_delay_1_payload_stateElements_9 <= partialRound_tempInput_payload_stateElements_9;
    partialRound_tempInput_delay_1_payload_stateElements_10 <= partialRound_tempInput_payload_stateElements_10;
    partialRound_tempInput_delay_1_payload_stateElements_11 <= partialRound_tempInput_payload_stateElements_11;
    partialRound_tempInput_delay_2_valid <= partialRound_tempInput_delay_1_valid;
    partialRound_tempInput_delay_2_payload_isFull <= partialRound_tempInput_delay_1_payload_isFull;
    partialRound_tempInput_delay_2_payload_fullRound <= partialRound_tempInput_delay_1_payload_fullRound;
    partialRound_tempInput_delay_2_payload_partialRound <= partialRound_tempInput_delay_1_payload_partialRound;
    partialRound_tempInput_delay_2_payload_stateSize <= partialRound_tempInput_delay_1_payload_stateSize;
    partialRound_tempInput_delay_2_payload_stateID <= partialRound_tempInput_delay_1_payload_stateID;
    partialRound_tempInput_delay_2_payload_stateElements_0 <= partialRound_tempInput_delay_1_payload_stateElements_0;
    partialRound_tempInput_delay_2_payload_stateElements_1 <= partialRound_tempInput_delay_1_payload_stateElements_1;
    partialRound_tempInput_delay_2_payload_stateElements_2 <= partialRound_tempInput_delay_1_payload_stateElements_2;
    partialRound_tempInput_delay_2_payload_stateElements_3 <= partialRound_tempInput_delay_1_payload_stateElements_3;
    partialRound_tempInput_delay_2_payload_stateElements_4 <= partialRound_tempInput_delay_1_payload_stateElements_4;
    partialRound_tempInput_delay_2_payload_stateElements_5 <= partialRound_tempInput_delay_1_payload_stateElements_5;
    partialRound_tempInput_delay_2_payload_stateElements_6 <= partialRound_tempInput_delay_1_payload_stateElements_6;
    partialRound_tempInput_delay_2_payload_stateElements_7 <= partialRound_tempInput_delay_1_payload_stateElements_7;
    partialRound_tempInput_delay_2_payload_stateElements_8 <= partialRound_tempInput_delay_1_payload_stateElements_8;
    partialRound_tempInput_delay_2_payload_stateElements_9 <= partialRound_tempInput_delay_1_payload_stateElements_9;
    partialRound_tempInput_delay_2_payload_stateElements_10 <= partialRound_tempInput_delay_1_payload_stateElements_10;
    partialRound_tempInput_delay_2_payload_stateElements_11 <= partialRound_tempInput_delay_1_payload_stateElements_11;
    partialRound_tempInput_delay_3_valid <= partialRound_tempInput_delay_2_valid;
    partialRound_tempInput_delay_3_payload_isFull <= partialRound_tempInput_delay_2_payload_isFull;
    partialRound_tempInput_delay_3_payload_fullRound <= partialRound_tempInput_delay_2_payload_fullRound;
    partialRound_tempInput_delay_3_payload_partialRound <= partialRound_tempInput_delay_2_payload_partialRound;
    partialRound_tempInput_delay_3_payload_stateSize <= partialRound_tempInput_delay_2_payload_stateSize;
    partialRound_tempInput_delay_3_payload_stateID <= partialRound_tempInput_delay_2_payload_stateID;
    partialRound_tempInput_delay_3_payload_stateElements_0 <= partialRound_tempInput_delay_2_payload_stateElements_0;
    partialRound_tempInput_delay_3_payload_stateElements_1 <= partialRound_tempInput_delay_2_payload_stateElements_1;
    partialRound_tempInput_delay_3_payload_stateElements_2 <= partialRound_tempInput_delay_2_payload_stateElements_2;
    partialRound_tempInput_delay_3_payload_stateElements_3 <= partialRound_tempInput_delay_2_payload_stateElements_3;
    partialRound_tempInput_delay_3_payload_stateElements_4 <= partialRound_tempInput_delay_2_payload_stateElements_4;
    partialRound_tempInput_delay_3_payload_stateElements_5 <= partialRound_tempInput_delay_2_payload_stateElements_5;
    partialRound_tempInput_delay_3_payload_stateElements_6 <= partialRound_tempInput_delay_2_payload_stateElements_6;
    partialRound_tempInput_delay_3_payload_stateElements_7 <= partialRound_tempInput_delay_2_payload_stateElements_7;
    partialRound_tempInput_delay_3_payload_stateElements_8 <= partialRound_tempInput_delay_2_payload_stateElements_8;
    partialRound_tempInput_delay_3_payload_stateElements_9 <= partialRound_tempInput_delay_2_payload_stateElements_9;
    partialRound_tempInput_delay_3_payload_stateElements_10 <= partialRound_tempInput_delay_2_payload_stateElements_10;
    partialRound_tempInput_delay_3_payload_stateElements_11 <= partialRound_tempInput_delay_2_payload_stateElements_11;
    partialRound_tempInput_delay_4_valid <= partialRound_tempInput_delay_3_valid;
    partialRound_tempInput_delay_4_payload_isFull <= partialRound_tempInput_delay_3_payload_isFull;
    partialRound_tempInput_delay_4_payload_fullRound <= partialRound_tempInput_delay_3_payload_fullRound;
    partialRound_tempInput_delay_4_payload_partialRound <= partialRound_tempInput_delay_3_payload_partialRound;
    partialRound_tempInput_delay_4_payload_stateSize <= partialRound_tempInput_delay_3_payload_stateSize;
    partialRound_tempInput_delay_4_payload_stateID <= partialRound_tempInput_delay_3_payload_stateID;
    partialRound_tempInput_delay_4_payload_stateElements_0 <= partialRound_tempInput_delay_3_payload_stateElements_0;
    partialRound_tempInput_delay_4_payload_stateElements_1 <= partialRound_tempInput_delay_3_payload_stateElements_1;
    partialRound_tempInput_delay_4_payload_stateElements_2 <= partialRound_tempInput_delay_3_payload_stateElements_2;
    partialRound_tempInput_delay_4_payload_stateElements_3 <= partialRound_tempInput_delay_3_payload_stateElements_3;
    partialRound_tempInput_delay_4_payload_stateElements_4 <= partialRound_tempInput_delay_3_payload_stateElements_4;
    partialRound_tempInput_delay_4_payload_stateElements_5 <= partialRound_tempInput_delay_3_payload_stateElements_5;
    partialRound_tempInput_delay_4_payload_stateElements_6 <= partialRound_tempInput_delay_3_payload_stateElements_6;
    partialRound_tempInput_delay_4_payload_stateElements_7 <= partialRound_tempInput_delay_3_payload_stateElements_7;
    partialRound_tempInput_delay_4_payload_stateElements_8 <= partialRound_tempInput_delay_3_payload_stateElements_8;
    partialRound_tempInput_delay_4_payload_stateElements_9 <= partialRound_tempInput_delay_3_payload_stateElements_9;
    partialRound_tempInput_delay_4_payload_stateElements_10 <= partialRound_tempInput_delay_3_payload_stateElements_10;
    partialRound_tempInput_delay_4_payload_stateElements_11 <= partialRound_tempInput_delay_3_payload_stateElements_11;
    partialRound_tempInput_delay_5_valid <= partialRound_tempInput_delay_4_valid;
    partialRound_tempInput_delay_5_payload_isFull <= partialRound_tempInput_delay_4_payload_isFull;
    partialRound_tempInput_delay_5_payload_fullRound <= partialRound_tempInput_delay_4_payload_fullRound;
    partialRound_tempInput_delay_5_payload_partialRound <= partialRound_tempInput_delay_4_payload_partialRound;
    partialRound_tempInput_delay_5_payload_stateSize <= partialRound_tempInput_delay_4_payload_stateSize;
    partialRound_tempInput_delay_5_payload_stateID <= partialRound_tempInput_delay_4_payload_stateID;
    partialRound_tempInput_delay_5_payload_stateElements_0 <= partialRound_tempInput_delay_4_payload_stateElements_0;
    partialRound_tempInput_delay_5_payload_stateElements_1 <= partialRound_tempInput_delay_4_payload_stateElements_1;
    partialRound_tempInput_delay_5_payload_stateElements_2 <= partialRound_tempInput_delay_4_payload_stateElements_2;
    partialRound_tempInput_delay_5_payload_stateElements_3 <= partialRound_tempInput_delay_4_payload_stateElements_3;
    partialRound_tempInput_delay_5_payload_stateElements_4 <= partialRound_tempInput_delay_4_payload_stateElements_4;
    partialRound_tempInput_delay_5_payload_stateElements_5 <= partialRound_tempInput_delay_4_payload_stateElements_5;
    partialRound_tempInput_delay_5_payload_stateElements_6 <= partialRound_tempInput_delay_4_payload_stateElements_6;
    partialRound_tempInput_delay_5_payload_stateElements_7 <= partialRound_tempInput_delay_4_payload_stateElements_7;
    partialRound_tempInput_delay_5_payload_stateElements_8 <= partialRound_tempInput_delay_4_payload_stateElements_8;
    partialRound_tempInput_delay_5_payload_stateElements_9 <= partialRound_tempInput_delay_4_payload_stateElements_9;
    partialRound_tempInput_delay_5_payload_stateElements_10 <= partialRound_tempInput_delay_4_payload_stateElements_10;
    partialRound_tempInput_delay_5_payload_stateElements_11 <= partialRound_tempInput_delay_4_payload_stateElements_11;
    partialRound_tempInput_delay_6_valid <= partialRound_tempInput_delay_5_valid;
    partialRound_tempInput_delay_6_payload_isFull <= partialRound_tempInput_delay_5_payload_isFull;
    partialRound_tempInput_delay_6_payload_fullRound <= partialRound_tempInput_delay_5_payload_fullRound;
    partialRound_tempInput_delay_6_payload_partialRound <= partialRound_tempInput_delay_5_payload_partialRound;
    partialRound_tempInput_delay_6_payload_stateSize <= partialRound_tempInput_delay_5_payload_stateSize;
    partialRound_tempInput_delay_6_payload_stateID <= partialRound_tempInput_delay_5_payload_stateID;
    partialRound_tempInput_delay_6_payload_stateElements_0 <= partialRound_tempInput_delay_5_payload_stateElements_0;
    partialRound_tempInput_delay_6_payload_stateElements_1 <= partialRound_tempInput_delay_5_payload_stateElements_1;
    partialRound_tempInput_delay_6_payload_stateElements_2 <= partialRound_tempInput_delay_5_payload_stateElements_2;
    partialRound_tempInput_delay_6_payload_stateElements_3 <= partialRound_tempInput_delay_5_payload_stateElements_3;
    partialRound_tempInput_delay_6_payload_stateElements_4 <= partialRound_tempInput_delay_5_payload_stateElements_4;
    partialRound_tempInput_delay_6_payload_stateElements_5 <= partialRound_tempInput_delay_5_payload_stateElements_5;
    partialRound_tempInput_delay_6_payload_stateElements_6 <= partialRound_tempInput_delay_5_payload_stateElements_6;
    partialRound_tempInput_delay_6_payload_stateElements_7 <= partialRound_tempInput_delay_5_payload_stateElements_7;
    partialRound_tempInput_delay_6_payload_stateElements_8 <= partialRound_tempInput_delay_5_payload_stateElements_8;
    partialRound_tempInput_delay_6_payload_stateElements_9 <= partialRound_tempInput_delay_5_payload_stateElements_9;
    partialRound_tempInput_delay_6_payload_stateElements_10 <= partialRound_tempInput_delay_5_payload_stateElements_10;
    partialRound_tempInput_delay_6_payload_stateElements_11 <= partialRound_tempInput_delay_5_payload_stateElements_11;
    partialRound_tempInput_delay_7_valid <= partialRound_tempInput_delay_6_valid;
    partialRound_tempInput_delay_7_payload_isFull <= partialRound_tempInput_delay_6_payload_isFull;
    partialRound_tempInput_delay_7_payload_fullRound <= partialRound_tempInput_delay_6_payload_fullRound;
    partialRound_tempInput_delay_7_payload_partialRound <= partialRound_tempInput_delay_6_payload_partialRound;
    partialRound_tempInput_delay_7_payload_stateSize <= partialRound_tempInput_delay_6_payload_stateSize;
    partialRound_tempInput_delay_7_payload_stateID <= partialRound_tempInput_delay_6_payload_stateID;
    partialRound_tempInput_delay_7_payload_stateElements_0 <= partialRound_tempInput_delay_6_payload_stateElements_0;
    partialRound_tempInput_delay_7_payload_stateElements_1 <= partialRound_tempInput_delay_6_payload_stateElements_1;
    partialRound_tempInput_delay_7_payload_stateElements_2 <= partialRound_tempInput_delay_6_payload_stateElements_2;
    partialRound_tempInput_delay_7_payload_stateElements_3 <= partialRound_tempInput_delay_6_payload_stateElements_3;
    partialRound_tempInput_delay_7_payload_stateElements_4 <= partialRound_tempInput_delay_6_payload_stateElements_4;
    partialRound_tempInput_delay_7_payload_stateElements_5 <= partialRound_tempInput_delay_6_payload_stateElements_5;
    partialRound_tempInput_delay_7_payload_stateElements_6 <= partialRound_tempInput_delay_6_payload_stateElements_6;
    partialRound_tempInput_delay_7_payload_stateElements_7 <= partialRound_tempInput_delay_6_payload_stateElements_7;
    partialRound_tempInput_delay_7_payload_stateElements_8 <= partialRound_tempInput_delay_6_payload_stateElements_8;
    partialRound_tempInput_delay_7_payload_stateElements_9 <= partialRound_tempInput_delay_6_payload_stateElements_9;
    partialRound_tempInput_delay_7_payload_stateElements_10 <= partialRound_tempInput_delay_6_payload_stateElements_10;
    partialRound_tempInput_delay_7_payload_stateElements_11 <= partialRound_tempInput_delay_6_payload_stateElements_11;
    partialRound_tempInput_delay_8_valid <= partialRound_tempInput_delay_7_valid;
    partialRound_tempInput_delay_8_payload_isFull <= partialRound_tempInput_delay_7_payload_isFull;
    partialRound_tempInput_delay_8_payload_fullRound <= partialRound_tempInput_delay_7_payload_fullRound;
    partialRound_tempInput_delay_8_payload_partialRound <= partialRound_tempInput_delay_7_payload_partialRound;
    partialRound_tempInput_delay_8_payload_stateSize <= partialRound_tempInput_delay_7_payload_stateSize;
    partialRound_tempInput_delay_8_payload_stateID <= partialRound_tempInput_delay_7_payload_stateID;
    partialRound_tempInput_delay_8_payload_stateElements_0 <= partialRound_tempInput_delay_7_payload_stateElements_0;
    partialRound_tempInput_delay_8_payload_stateElements_1 <= partialRound_tempInput_delay_7_payload_stateElements_1;
    partialRound_tempInput_delay_8_payload_stateElements_2 <= partialRound_tempInput_delay_7_payload_stateElements_2;
    partialRound_tempInput_delay_8_payload_stateElements_3 <= partialRound_tempInput_delay_7_payload_stateElements_3;
    partialRound_tempInput_delay_8_payload_stateElements_4 <= partialRound_tempInput_delay_7_payload_stateElements_4;
    partialRound_tempInput_delay_8_payload_stateElements_5 <= partialRound_tempInput_delay_7_payload_stateElements_5;
    partialRound_tempInput_delay_8_payload_stateElements_6 <= partialRound_tempInput_delay_7_payload_stateElements_6;
    partialRound_tempInput_delay_8_payload_stateElements_7 <= partialRound_tempInput_delay_7_payload_stateElements_7;
    partialRound_tempInput_delay_8_payload_stateElements_8 <= partialRound_tempInput_delay_7_payload_stateElements_8;
    partialRound_tempInput_delay_8_payload_stateElements_9 <= partialRound_tempInput_delay_7_payload_stateElements_9;
    partialRound_tempInput_delay_8_payload_stateElements_10 <= partialRound_tempInput_delay_7_payload_stateElements_10;
    partialRound_tempInput_delay_8_payload_stateElements_11 <= partialRound_tempInput_delay_7_payload_stateElements_11;
    partialRound_tempInput_delay_9_valid <= partialRound_tempInput_delay_8_valid;
    partialRound_tempInput_delay_9_payload_isFull <= partialRound_tempInput_delay_8_payload_isFull;
    partialRound_tempInput_delay_9_payload_fullRound <= partialRound_tempInput_delay_8_payload_fullRound;
    partialRound_tempInput_delay_9_payload_partialRound <= partialRound_tempInput_delay_8_payload_partialRound;
    partialRound_tempInput_delay_9_payload_stateSize <= partialRound_tempInput_delay_8_payload_stateSize;
    partialRound_tempInput_delay_9_payload_stateID <= partialRound_tempInput_delay_8_payload_stateID;
    partialRound_tempInput_delay_9_payload_stateElements_0 <= partialRound_tempInput_delay_8_payload_stateElements_0;
    partialRound_tempInput_delay_9_payload_stateElements_1 <= partialRound_tempInput_delay_8_payload_stateElements_1;
    partialRound_tempInput_delay_9_payload_stateElements_2 <= partialRound_tempInput_delay_8_payload_stateElements_2;
    partialRound_tempInput_delay_9_payload_stateElements_3 <= partialRound_tempInput_delay_8_payload_stateElements_3;
    partialRound_tempInput_delay_9_payload_stateElements_4 <= partialRound_tempInput_delay_8_payload_stateElements_4;
    partialRound_tempInput_delay_9_payload_stateElements_5 <= partialRound_tempInput_delay_8_payload_stateElements_5;
    partialRound_tempInput_delay_9_payload_stateElements_6 <= partialRound_tempInput_delay_8_payload_stateElements_6;
    partialRound_tempInput_delay_9_payload_stateElements_7 <= partialRound_tempInput_delay_8_payload_stateElements_7;
    partialRound_tempInput_delay_9_payload_stateElements_8 <= partialRound_tempInput_delay_8_payload_stateElements_8;
    partialRound_tempInput_delay_9_payload_stateElements_9 <= partialRound_tempInput_delay_8_payload_stateElements_9;
    partialRound_tempInput_delay_9_payload_stateElements_10 <= partialRound_tempInput_delay_8_payload_stateElements_10;
    partialRound_tempInput_delay_9_payload_stateElements_11 <= partialRound_tempInput_delay_8_payload_stateElements_11;
    partialRound_tempInput_delay_10_valid <= partialRound_tempInput_delay_9_valid;
    partialRound_tempInput_delay_10_payload_isFull <= partialRound_tempInput_delay_9_payload_isFull;
    partialRound_tempInput_delay_10_payload_fullRound <= partialRound_tempInput_delay_9_payload_fullRound;
    partialRound_tempInput_delay_10_payload_partialRound <= partialRound_tempInput_delay_9_payload_partialRound;
    partialRound_tempInput_delay_10_payload_stateSize <= partialRound_tempInput_delay_9_payload_stateSize;
    partialRound_tempInput_delay_10_payload_stateID <= partialRound_tempInput_delay_9_payload_stateID;
    partialRound_tempInput_delay_10_payload_stateElements_0 <= partialRound_tempInput_delay_9_payload_stateElements_0;
    partialRound_tempInput_delay_10_payload_stateElements_1 <= partialRound_tempInput_delay_9_payload_stateElements_1;
    partialRound_tempInput_delay_10_payload_stateElements_2 <= partialRound_tempInput_delay_9_payload_stateElements_2;
    partialRound_tempInput_delay_10_payload_stateElements_3 <= partialRound_tempInput_delay_9_payload_stateElements_3;
    partialRound_tempInput_delay_10_payload_stateElements_4 <= partialRound_tempInput_delay_9_payload_stateElements_4;
    partialRound_tempInput_delay_10_payload_stateElements_5 <= partialRound_tempInput_delay_9_payload_stateElements_5;
    partialRound_tempInput_delay_10_payload_stateElements_6 <= partialRound_tempInput_delay_9_payload_stateElements_6;
    partialRound_tempInput_delay_10_payload_stateElements_7 <= partialRound_tempInput_delay_9_payload_stateElements_7;
    partialRound_tempInput_delay_10_payload_stateElements_8 <= partialRound_tempInput_delay_9_payload_stateElements_8;
    partialRound_tempInput_delay_10_payload_stateElements_9 <= partialRound_tempInput_delay_9_payload_stateElements_9;
    partialRound_tempInput_delay_10_payload_stateElements_10 <= partialRound_tempInput_delay_9_payload_stateElements_10;
    partialRound_tempInput_delay_10_payload_stateElements_11 <= partialRound_tempInput_delay_9_payload_stateElements_11;
    partialRound_tempInput_delay_11_valid <= partialRound_tempInput_delay_10_valid;
    partialRound_tempInput_delay_11_payload_isFull <= partialRound_tempInput_delay_10_payload_isFull;
    partialRound_tempInput_delay_11_payload_fullRound <= partialRound_tempInput_delay_10_payload_fullRound;
    partialRound_tempInput_delay_11_payload_partialRound <= partialRound_tempInput_delay_10_payload_partialRound;
    partialRound_tempInput_delay_11_payload_stateSize <= partialRound_tempInput_delay_10_payload_stateSize;
    partialRound_tempInput_delay_11_payload_stateID <= partialRound_tempInput_delay_10_payload_stateID;
    partialRound_tempInput_delay_11_payload_stateElements_0 <= partialRound_tempInput_delay_10_payload_stateElements_0;
    partialRound_tempInput_delay_11_payload_stateElements_1 <= partialRound_tempInput_delay_10_payload_stateElements_1;
    partialRound_tempInput_delay_11_payload_stateElements_2 <= partialRound_tempInput_delay_10_payload_stateElements_2;
    partialRound_tempInput_delay_11_payload_stateElements_3 <= partialRound_tempInput_delay_10_payload_stateElements_3;
    partialRound_tempInput_delay_11_payload_stateElements_4 <= partialRound_tempInput_delay_10_payload_stateElements_4;
    partialRound_tempInput_delay_11_payload_stateElements_5 <= partialRound_tempInput_delay_10_payload_stateElements_5;
    partialRound_tempInput_delay_11_payload_stateElements_6 <= partialRound_tempInput_delay_10_payload_stateElements_6;
    partialRound_tempInput_delay_11_payload_stateElements_7 <= partialRound_tempInput_delay_10_payload_stateElements_7;
    partialRound_tempInput_delay_11_payload_stateElements_8 <= partialRound_tempInput_delay_10_payload_stateElements_8;
    partialRound_tempInput_delay_11_payload_stateElements_9 <= partialRound_tempInput_delay_10_payload_stateElements_9;
    partialRound_tempInput_delay_11_payload_stateElements_10 <= partialRound_tempInput_delay_10_payload_stateElements_10;
    partialRound_tempInput_delay_11_payload_stateElements_11 <= partialRound_tempInput_delay_10_payload_stateElements_11;
    partialRound_tempInput_delay_12_valid <= partialRound_tempInput_delay_11_valid;
    partialRound_tempInput_delay_12_payload_isFull <= partialRound_tempInput_delay_11_payload_isFull;
    partialRound_tempInput_delay_12_payload_fullRound <= partialRound_tempInput_delay_11_payload_fullRound;
    partialRound_tempInput_delay_12_payload_partialRound <= partialRound_tempInput_delay_11_payload_partialRound;
    partialRound_tempInput_delay_12_payload_stateSize <= partialRound_tempInput_delay_11_payload_stateSize;
    partialRound_tempInput_delay_12_payload_stateID <= partialRound_tempInput_delay_11_payload_stateID;
    partialRound_tempInput_delay_12_payload_stateElements_0 <= partialRound_tempInput_delay_11_payload_stateElements_0;
    partialRound_tempInput_delay_12_payload_stateElements_1 <= partialRound_tempInput_delay_11_payload_stateElements_1;
    partialRound_tempInput_delay_12_payload_stateElements_2 <= partialRound_tempInput_delay_11_payload_stateElements_2;
    partialRound_tempInput_delay_12_payload_stateElements_3 <= partialRound_tempInput_delay_11_payload_stateElements_3;
    partialRound_tempInput_delay_12_payload_stateElements_4 <= partialRound_tempInput_delay_11_payload_stateElements_4;
    partialRound_tempInput_delay_12_payload_stateElements_5 <= partialRound_tempInput_delay_11_payload_stateElements_5;
    partialRound_tempInput_delay_12_payload_stateElements_6 <= partialRound_tempInput_delay_11_payload_stateElements_6;
    partialRound_tempInput_delay_12_payload_stateElements_7 <= partialRound_tempInput_delay_11_payload_stateElements_7;
    partialRound_tempInput_delay_12_payload_stateElements_8 <= partialRound_tempInput_delay_11_payload_stateElements_8;
    partialRound_tempInput_delay_12_payload_stateElements_9 <= partialRound_tempInput_delay_11_payload_stateElements_9;
    partialRound_tempInput_delay_12_payload_stateElements_10 <= partialRound_tempInput_delay_11_payload_stateElements_10;
    partialRound_tempInput_delay_12_payload_stateElements_11 <= partialRound_tempInput_delay_11_payload_stateElements_11;
    partialRound_tempInput_delay_13_valid <= partialRound_tempInput_delay_12_valid;
    partialRound_tempInput_delay_13_payload_isFull <= partialRound_tempInput_delay_12_payload_isFull;
    partialRound_tempInput_delay_13_payload_fullRound <= partialRound_tempInput_delay_12_payload_fullRound;
    partialRound_tempInput_delay_13_payload_partialRound <= partialRound_tempInput_delay_12_payload_partialRound;
    partialRound_tempInput_delay_13_payload_stateSize <= partialRound_tempInput_delay_12_payload_stateSize;
    partialRound_tempInput_delay_13_payload_stateID <= partialRound_tempInput_delay_12_payload_stateID;
    partialRound_tempInput_delay_13_payload_stateElements_0 <= partialRound_tempInput_delay_12_payload_stateElements_0;
    partialRound_tempInput_delay_13_payload_stateElements_1 <= partialRound_tempInput_delay_12_payload_stateElements_1;
    partialRound_tempInput_delay_13_payload_stateElements_2 <= partialRound_tempInput_delay_12_payload_stateElements_2;
    partialRound_tempInput_delay_13_payload_stateElements_3 <= partialRound_tempInput_delay_12_payload_stateElements_3;
    partialRound_tempInput_delay_13_payload_stateElements_4 <= partialRound_tempInput_delay_12_payload_stateElements_4;
    partialRound_tempInput_delay_13_payload_stateElements_5 <= partialRound_tempInput_delay_12_payload_stateElements_5;
    partialRound_tempInput_delay_13_payload_stateElements_6 <= partialRound_tempInput_delay_12_payload_stateElements_6;
    partialRound_tempInput_delay_13_payload_stateElements_7 <= partialRound_tempInput_delay_12_payload_stateElements_7;
    partialRound_tempInput_delay_13_payload_stateElements_8 <= partialRound_tempInput_delay_12_payload_stateElements_8;
    partialRound_tempInput_delay_13_payload_stateElements_9 <= partialRound_tempInput_delay_12_payload_stateElements_9;
    partialRound_tempInput_delay_13_payload_stateElements_10 <= partialRound_tempInput_delay_12_payload_stateElements_10;
    partialRound_tempInput_delay_13_payload_stateElements_11 <= partialRound_tempInput_delay_12_payload_stateElements_11;
    partialRound_tempInput_delay_14_valid <= partialRound_tempInput_delay_13_valid;
    partialRound_tempInput_delay_14_payload_isFull <= partialRound_tempInput_delay_13_payload_isFull;
    partialRound_tempInput_delay_14_payload_fullRound <= partialRound_tempInput_delay_13_payload_fullRound;
    partialRound_tempInput_delay_14_payload_partialRound <= partialRound_tempInput_delay_13_payload_partialRound;
    partialRound_tempInput_delay_14_payload_stateSize <= partialRound_tempInput_delay_13_payload_stateSize;
    partialRound_tempInput_delay_14_payload_stateID <= partialRound_tempInput_delay_13_payload_stateID;
    partialRound_tempInput_delay_14_payload_stateElements_0 <= partialRound_tempInput_delay_13_payload_stateElements_0;
    partialRound_tempInput_delay_14_payload_stateElements_1 <= partialRound_tempInput_delay_13_payload_stateElements_1;
    partialRound_tempInput_delay_14_payload_stateElements_2 <= partialRound_tempInput_delay_13_payload_stateElements_2;
    partialRound_tempInput_delay_14_payload_stateElements_3 <= partialRound_tempInput_delay_13_payload_stateElements_3;
    partialRound_tempInput_delay_14_payload_stateElements_4 <= partialRound_tempInput_delay_13_payload_stateElements_4;
    partialRound_tempInput_delay_14_payload_stateElements_5 <= partialRound_tempInput_delay_13_payload_stateElements_5;
    partialRound_tempInput_delay_14_payload_stateElements_6 <= partialRound_tempInput_delay_13_payload_stateElements_6;
    partialRound_tempInput_delay_14_payload_stateElements_7 <= partialRound_tempInput_delay_13_payload_stateElements_7;
    partialRound_tempInput_delay_14_payload_stateElements_8 <= partialRound_tempInput_delay_13_payload_stateElements_8;
    partialRound_tempInput_delay_14_payload_stateElements_9 <= partialRound_tempInput_delay_13_payload_stateElements_9;
    partialRound_tempInput_delay_14_payload_stateElements_10 <= partialRound_tempInput_delay_13_payload_stateElements_10;
    partialRound_tempInput_delay_14_payload_stateElements_11 <= partialRound_tempInput_delay_13_payload_stateElements_11;
    partialRound_tempInput_delay_15_valid <= partialRound_tempInput_delay_14_valid;
    partialRound_tempInput_delay_15_payload_isFull <= partialRound_tempInput_delay_14_payload_isFull;
    partialRound_tempInput_delay_15_payload_fullRound <= partialRound_tempInput_delay_14_payload_fullRound;
    partialRound_tempInput_delay_15_payload_partialRound <= partialRound_tempInput_delay_14_payload_partialRound;
    partialRound_tempInput_delay_15_payload_stateSize <= partialRound_tempInput_delay_14_payload_stateSize;
    partialRound_tempInput_delay_15_payload_stateID <= partialRound_tempInput_delay_14_payload_stateID;
    partialRound_tempInput_delay_15_payload_stateElements_0 <= partialRound_tempInput_delay_14_payload_stateElements_0;
    partialRound_tempInput_delay_15_payload_stateElements_1 <= partialRound_tempInput_delay_14_payload_stateElements_1;
    partialRound_tempInput_delay_15_payload_stateElements_2 <= partialRound_tempInput_delay_14_payload_stateElements_2;
    partialRound_tempInput_delay_15_payload_stateElements_3 <= partialRound_tempInput_delay_14_payload_stateElements_3;
    partialRound_tempInput_delay_15_payload_stateElements_4 <= partialRound_tempInput_delay_14_payload_stateElements_4;
    partialRound_tempInput_delay_15_payload_stateElements_5 <= partialRound_tempInput_delay_14_payload_stateElements_5;
    partialRound_tempInput_delay_15_payload_stateElements_6 <= partialRound_tempInput_delay_14_payload_stateElements_6;
    partialRound_tempInput_delay_15_payload_stateElements_7 <= partialRound_tempInput_delay_14_payload_stateElements_7;
    partialRound_tempInput_delay_15_payload_stateElements_8 <= partialRound_tempInput_delay_14_payload_stateElements_8;
    partialRound_tempInput_delay_15_payload_stateElements_9 <= partialRound_tempInput_delay_14_payload_stateElements_9;
    partialRound_tempInput_delay_15_payload_stateElements_10 <= partialRound_tempInput_delay_14_payload_stateElements_10;
    partialRound_tempInput_delay_15_payload_stateElements_11 <= partialRound_tempInput_delay_14_payload_stateElements_11;
    partialRound_tempInput_delay_16_valid <= partialRound_tempInput_delay_15_valid;
    partialRound_tempInput_delay_16_payload_isFull <= partialRound_tempInput_delay_15_payload_isFull;
    partialRound_tempInput_delay_16_payload_fullRound <= partialRound_tempInput_delay_15_payload_fullRound;
    partialRound_tempInput_delay_16_payload_partialRound <= partialRound_tempInput_delay_15_payload_partialRound;
    partialRound_tempInput_delay_16_payload_stateSize <= partialRound_tempInput_delay_15_payload_stateSize;
    partialRound_tempInput_delay_16_payload_stateID <= partialRound_tempInput_delay_15_payload_stateID;
    partialRound_tempInput_delay_16_payload_stateElements_0 <= partialRound_tempInput_delay_15_payload_stateElements_0;
    partialRound_tempInput_delay_16_payload_stateElements_1 <= partialRound_tempInput_delay_15_payload_stateElements_1;
    partialRound_tempInput_delay_16_payload_stateElements_2 <= partialRound_tempInput_delay_15_payload_stateElements_2;
    partialRound_tempInput_delay_16_payload_stateElements_3 <= partialRound_tempInput_delay_15_payload_stateElements_3;
    partialRound_tempInput_delay_16_payload_stateElements_4 <= partialRound_tempInput_delay_15_payload_stateElements_4;
    partialRound_tempInput_delay_16_payload_stateElements_5 <= partialRound_tempInput_delay_15_payload_stateElements_5;
    partialRound_tempInput_delay_16_payload_stateElements_6 <= partialRound_tempInput_delay_15_payload_stateElements_6;
    partialRound_tempInput_delay_16_payload_stateElements_7 <= partialRound_tempInput_delay_15_payload_stateElements_7;
    partialRound_tempInput_delay_16_payload_stateElements_8 <= partialRound_tempInput_delay_15_payload_stateElements_8;
    partialRound_tempInput_delay_16_payload_stateElements_9 <= partialRound_tempInput_delay_15_payload_stateElements_9;
    partialRound_tempInput_delay_16_payload_stateElements_10 <= partialRound_tempInput_delay_15_payload_stateElements_10;
    partialRound_tempInput_delay_16_payload_stateElements_11 <= partialRound_tempInput_delay_15_payload_stateElements_11;
    partialRound_tempInput_delay_17_valid <= partialRound_tempInput_delay_16_valid;
    partialRound_tempInput_delay_17_payload_isFull <= partialRound_tempInput_delay_16_payload_isFull;
    partialRound_tempInput_delay_17_payload_fullRound <= partialRound_tempInput_delay_16_payload_fullRound;
    partialRound_tempInput_delay_17_payload_partialRound <= partialRound_tempInput_delay_16_payload_partialRound;
    partialRound_tempInput_delay_17_payload_stateSize <= partialRound_tempInput_delay_16_payload_stateSize;
    partialRound_tempInput_delay_17_payload_stateID <= partialRound_tempInput_delay_16_payload_stateID;
    partialRound_tempInput_delay_17_payload_stateElements_0 <= partialRound_tempInput_delay_16_payload_stateElements_0;
    partialRound_tempInput_delay_17_payload_stateElements_1 <= partialRound_tempInput_delay_16_payload_stateElements_1;
    partialRound_tempInput_delay_17_payload_stateElements_2 <= partialRound_tempInput_delay_16_payload_stateElements_2;
    partialRound_tempInput_delay_17_payload_stateElements_3 <= partialRound_tempInput_delay_16_payload_stateElements_3;
    partialRound_tempInput_delay_17_payload_stateElements_4 <= partialRound_tempInput_delay_16_payload_stateElements_4;
    partialRound_tempInput_delay_17_payload_stateElements_5 <= partialRound_tempInput_delay_16_payload_stateElements_5;
    partialRound_tempInput_delay_17_payload_stateElements_6 <= partialRound_tempInput_delay_16_payload_stateElements_6;
    partialRound_tempInput_delay_17_payload_stateElements_7 <= partialRound_tempInput_delay_16_payload_stateElements_7;
    partialRound_tempInput_delay_17_payload_stateElements_8 <= partialRound_tempInput_delay_16_payload_stateElements_8;
    partialRound_tempInput_delay_17_payload_stateElements_9 <= partialRound_tempInput_delay_16_payload_stateElements_9;
    partialRound_tempInput_delay_17_payload_stateElements_10 <= partialRound_tempInput_delay_16_payload_stateElements_10;
    partialRound_tempInput_delay_17_payload_stateElements_11 <= partialRound_tempInput_delay_16_payload_stateElements_11;
    partialRound_tempInput_delay_18_valid <= partialRound_tempInput_delay_17_valid;
    partialRound_tempInput_delay_18_payload_isFull <= partialRound_tempInput_delay_17_payload_isFull;
    partialRound_tempInput_delay_18_payload_fullRound <= partialRound_tempInput_delay_17_payload_fullRound;
    partialRound_tempInput_delay_18_payload_partialRound <= partialRound_tempInput_delay_17_payload_partialRound;
    partialRound_tempInput_delay_18_payload_stateSize <= partialRound_tempInput_delay_17_payload_stateSize;
    partialRound_tempInput_delay_18_payload_stateID <= partialRound_tempInput_delay_17_payload_stateID;
    partialRound_tempInput_delay_18_payload_stateElements_0 <= partialRound_tempInput_delay_17_payload_stateElements_0;
    partialRound_tempInput_delay_18_payload_stateElements_1 <= partialRound_tempInput_delay_17_payload_stateElements_1;
    partialRound_tempInput_delay_18_payload_stateElements_2 <= partialRound_tempInput_delay_17_payload_stateElements_2;
    partialRound_tempInput_delay_18_payload_stateElements_3 <= partialRound_tempInput_delay_17_payload_stateElements_3;
    partialRound_tempInput_delay_18_payload_stateElements_4 <= partialRound_tempInput_delay_17_payload_stateElements_4;
    partialRound_tempInput_delay_18_payload_stateElements_5 <= partialRound_tempInput_delay_17_payload_stateElements_5;
    partialRound_tempInput_delay_18_payload_stateElements_6 <= partialRound_tempInput_delay_17_payload_stateElements_6;
    partialRound_tempInput_delay_18_payload_stateElements_7 <= partialRound_tempInput_delay_17_payload_stateElements_7;
    partialRound_tempInput_delay_18_payload_stateElements_8 <= partialRound_tempInput_delay_17_payload_stateElements_8;
    partialRound_tempInput_delay_18_payload_stateElements_9 <= partialRound_tempInput_delay_17_payload_stateElements_9;
    partialRound_tempInput_delay_18_payload_stateElements_10 <= partialRound_tempInput_delay_17_payload_stateElements_10;
    partialRound_tempInput_delay_18_payload_stateElements_11 <= partialRound_tempInput_delay_17_payload_stateElements_11;
    partialRound_tempInput_delay_19_valid <= partialRound_tempInput_delay_18_valid;
    partialRound_tempInput_delay_19_payload_isFull <= partialRound_tempInput_delay_18_payload_isFull;
    partialRound_tempInput_delay_19_payload_fullRound <= partialRound_tempInput_delay_18_payload_fullRound;
    partialRound_tempInput_delay_19_payload_partialRound <= partialRound_tempInput_delay_18_payload_partialRound;
    partialRound_tempInput_delay_19_payload_stateSize <= partialRound_tempInput_delay_18_payload_stateSize;
    partialRound_tempInput_delay_19_payload_stateID <= partialRound_tempInput_delay_18_payload_stateID;
    partialRound_tempInput_delay_19_payload_stateElements_0 <= partialRound_tempInput_delay_18_payload_stateElements_0;
    partialRound_tempInput_delay_19_payload_stateElements_1 <= partialRound_tempInput_delay_18_payload_stateElements_1;
    partialRound_tempInput_delay_19_payload_stateElements_2 <= partialRound_tempInput_delay_18_payload_stateElements_2;
    partialRound_tempInput_delay_19_payload_stateElements_3 <= partialRound_tempInput_delay_18_payload_stateElements_3;
    partialRound_tempInput_delay_19_payload_stateElements_4 <= partialRound_tempInput_delay_18_payload_stateElements_4;
    partialRound_tempInput_delay_19_payload_stateElements_5 <= partialRound_tempInput_delay_18_payload_stateElements_5;
    partialRound_tempInput_delay_19_payload_stateElements_6 <= partialRound_tempInput_delay_18_payload_stateElements_6;
    partialRound_tempInput_delay_19_payload_stateElements_7 <= partialRound_tempInput_delay_18_payload_stateElements_7;
    partialRound_tempInput_delay_19_payload_stateElements_8 <= partialRound_tempInput_delay_18_payload_stateElements_8;
    partialRound_tempInput_delay_19_payload_stateElements_9 <= partialRound_tempInput_delay_18_payload_stateElements_9;
    partialRound_tempInput_delay_19_payload_stateElements_10 <= partialRound_tempInput_delay_18_payload_stateElements_10;
    partialRound_tempInput_delay_19_payload_stateElements_11 <= partialRound_tempInput_delay_18_payload_stateElements_11;
    partialRound_tempInput_delay_20_valid <= partialRound_tempInput_delay_19_valid;
    partialRound_tempInput_delay_20_payload_isFull <= partialRound_tempInput_delay_19_payload_isFull;
    partialRound_tempInput_delay_20_payload_fullRound <= partialRound_tempInput_delay_19_payload_fullRound;
    partialRound_tempInput_delay_20_payload_partialRound <= partialRound_tempInput_delay_19_payload_partialRound;
    partialRound_tempInput_delay_20_payload_stateSize <= partialRound_tempInput_delay_19_payload_stateSize;
    partialRound_tempInput_delay_20_payload_stateID <= partialRound_tempInput_delay_19_payload_stateID;
    partialRound_tempInput_delay_20_payload_stateElements_0 <= partialRound_tempInput_delay_19_payload_stateElements_0;
    partialRound_tempInput_delay_20_payload_stateElements_1 <= partialRound_tempInput_delay_19_payload_stateElements_1;
    partialRound_tempInput_delay_20_payload_stateElements_2 <= partialRound_tempInput_delay_19_payload_stateElements_2;
    partialRound_tempInput_delay_20_payload_stateElements_3 <= partialRound_tempInput_delay_19_payload_stateElements_3;
    partialRound_tempInput_delay_20_payload_stateElements_4 <= partialRound_tempInput_delay_19_payload_stateElements_4;
    partialRound_tempInput_delay_20_payload_stateElements_5 <= partialRound_tempInput_delay_19_payload_stateElements_5;
    partialRound_tempInput_delay_20_payload_stateElements_6 <= partialRound_tempInput_delay_19_payload_stateElements_6;
    partialRound_tempInput_delay_20_payload_stateElements_7 <= partialRound_tempInput_delay_19_payload_stateElements_7;
    partialRound_tempInput_delay_20_payload_stateElements_8 <= partialRound_tempInput_delay_19_payload_stateElements_8;
    partialRound_tempInput_delay_20_payload_stateElements_9 <= partialRound_tempInput_delay_19_payload_stateElements_9;
    partialRound_tempInput_delay_20_payload_stateElements_10 <= partialRound_tempInput_delay_19_payload_stateElements_10;
    partialRound_tempInput_delay_20_payload_stateElements_11 <= partialRound_tempInput_delay_19_payload_stateElements_11;
    partialRound_tempInput_delay_21_valid <= partialRound_tempInput_delay_20_valid;
    partialRound_tempInput_delay_21_payload_isFull <= partialRound_tempInput_delay_20_payload_isFull;
    partialRound_tempInput_delay_21_payload_fullRound <= partialRound_tempInput_delay_20_payload_fullRound;
    partialRound_tempInput_delay_21_payload_partialRound <= partialRound_tempInput_delay_20_payload_partialRound;
    partialRound_tempInput_delay_21_payload_stateSize <= partialRound_tempInput_delay_20_payload_stateSize;
    partialRound_tempInput_delay_21_payload_stateID <= partialRound_tempInput_delay_20_payload_stateID;
    partialRound_tempInput_delay_21_payload_stateElements_0 <= partialRound_tempInput_delay_20_payload_stateElements_0;
    partialRound_tempInput_delay_21_payload_stateElements_1 <= partialRound_tempInput_delay_20_payload_stateElements_1;
    partialRound_tempInput_delay_21_payload_stateElements_2 <= partialRound_tempInput_delay_20_payload_stateElements_2;
    partialRound_tempInput_delay_21_payload_stateElements_3 <= partialRound_tempInput_delay_20_payload_stateElements_3;
    partialRound_tempInput_delay_21_payload_stateElements_4 <= partialRound_tempInput_delay_20_payload_stateElements_4;
    partialRound_tempInput_delay_21_payload_stateElements_5 <= partialRound_tempInput_delay_20_payload_stateElements_5;
    partialRound_tempInput_delay_21_payload_stateElements_6 <= partialRound_tempInput_delay_20_payload_stateElements_6;
    partialRound_tempInput_delay_21_payload_stateElements_7 <= partialRound_tempInput_delay_20_payload_stateElements_7;
    partialRound_tempInput_delay_21_payload_stateElements_8 <= partialRound_tempInput_delay_20_payload_stateElements_8;
    partialRound_tempInput_delay_21_payload_stateElements_9 <= partialRound_tempInput_delay_20_payload_stateElements_9;
    partialRound_tempInput_delay_21_payload_stateElements_10 <= partialRound_tempInput_delay_20_payload_stateElements_10;
    partialRound_tempInput_delay_21_payload_stateElements_11 <= partialRound_tempInput_delay_20_payload_stateElements_11;
    partialRound_tempInput_delay_22_valid <= partialRound_tempInput_delay_21_valid;
    partialRound_tempInput_delay_22_payload_isFull <= partialRound_tempInput_delay_21_payload_isFull;
    partialRound_tempInput_delay_22_payload_fullRound <= partialRound_tempInput_delay_21_payload_fullRound;
    partialRound_tempInput_delay_22_payload_partialRound <= partialRound_tempInput_delay_21_payload_partialRound;
    partialRound_tempInput_delay_22_payload_stateSize <= partialRound_tempInput_delay_21_payload_stateSize;
    partialRound_tempInput_delay_22_payload_stateID <= partialRound_tempInput_delay_21_payload_stateID;
    partialRound_tempInput_delay_22_payload_stateElements_0 <= partialRound_tempInput_delay_21_payload_stateElements_0;
    partialRound_tempInput_delay_22_payload_stateElements_1 <= partialRound_tempInput_delay_21_payload_stateElements_1;
    partialRound_tempInput_delay_22_payload_stateElements_2 <= partialRound_tempInput_delay_21_payload_stateElements_2;
    partialRound_tempInput_delay_22_payload_stateElements_3 <= partialRound_tempInput_delay_21_payload_stateElements_3;
    partialRound_tempInput_delay_22_payload_stateElements_4 <= partialRound_tempInput_delay_21_payload_stateElements_4;
    partialRound_tempInput_delay_22_payload_stateElements_5 <= partialRound_tempInput_delay_21_payload_stateElements_5;
    partialRound_tempInput_delay_22_payload_stateElements_6 <= partialRound_tempInput_delay_21_payload_stateElements_6;
    partialRound_tempInput_delay_22_payload_stateElements_7 <= partialRound_tempInput_delay_21_payload_stateElements_7;
    partialRound_tempInput_delay_22_payload_stateElements_8 <= partialRound_tempInput_delay_21_payload_stateElements_8;
    partialRound_tempInput_delay_22_payload_stateElements_9 <= partialRound_tempInput_delay_21_payload_stateElements_9;
    partialRound_tempInput_delay_22_payload_stateElements_10 <= partialRound_tempInput_delay_21_payload_stateElements_10;
    partialRound_tempInput_delay_22_payload_stateElements_11 <= partialRound_tempInput_delay_21_payload_stateElements_11;
    partialRound_tempInput_delay_23_valid <= partialRound_tempInput_delay_22_valid;
    partialRound_tempInput_delay_23_payload_isFull <= partialRound_tempInput_delay_22_payload_isFull;
    partialRound_tempInput_delay_23_payload_fullRound <= partialRound_tempInput_delay_22_payload_fullRound;
    partialRound_tempInput_delay_23_payload_partialRound <= partialRound_tempInput_delay_22_payload_partialRound;
    partialRound_tempInput_delay_23_payload_stateSize <= partialRound_tempInput_delay_22_payload_stateSize;
    partialRound_tempInput_delay_23_payload_stateID <= partialRound_tempInput_delay_22_payload_stateID;
    partialRound_tempInput_delay_23_payload_stateElements_0 <= partialRound_tempInput_delay_22_payload_stateElements_0;
    partialRound_tempInput_delay_23_payload_stateElements_1 <= partialRound_tempInput_delay_22_payload_stateElements_1;
    partialRound_tempInput_delay_23_payload_stateElements_2 <= partialRound_tempInput_delay_22_payload_stateElements_2;
    partialRound_tempInput_delay_23_payload_stateElements_3 <= partialRound_tempInput_delay_22_payload_stateElements_3;
    partialRound_tempInput_delay_23_payload_stateElements_4 <= partialRound_tempInput_delay_22_payload_stateElements_4;
    partialRound_tempInput_delay_23_payload_stateElements_5 <= partialRound_tempInput_delay_22_payload_stateElements_5;
    partialRound_tempInput_delay_23_payload_stateElements_6 <= partialRound_tempInput_delay_22_payload_stateElements_6;
    partialRound_tempInput_delay_23_payload_stateElements_7 <= partialRound_tempInput_delay_22_payload_stateElements_7;
    partialRound_tempInput_delay_23_payload_stateElements_8 <= partialRound_tempInput_delay_22_payload_stateElements_8;
    partialRound_tempInput_delay_23_payload_stateElements_9 <= partialRound_tempInput_delay_22_payload_stateElements_9;
    partialRound_tempInput_delay_23_payload_stateElements_10 <= partialRound_tempInput_delay_22_payload_stateElements_10;
    partialRound_tempInput_delay_23_payload_stateElements_11 <= partialRound_tempInput_delay_22_payload_stateElements_11;
    partialRound_tempInput_delay_24_valid <= partialRound_tempInput_delay_23_valid;
    partialRound_tempInput_delay_24_payload_isFull <= partialRound_tempInput_delay_23_payload_isFull;
    partialRound_tempInput_delay_24_payload_fullRound <= partialRound_tempInput_delay_23_payload_fullRound;
    partialRound_tempInput_delay_24_payload_partialRound <= partialRound_tempInput_delay_23_payload_partialRound;
    partialRound_tempInput_delay_24_payload_stateSize <= partialRound_tempInput_delay_23_payload_stateSize;
    partialRound_tempInput_delay_24_payload_stateID <= partialRound_tempInput_delay_23_payload_stateID;
    partialRound_tempInput_delay_24_payload_stateElements_0 <= partialRound_tempInput_delay_23_payload_stateElements_0;
    partialRound_tempInput_delay_24_payload_stateElements_1 <= partialRound_tempInput_delay_23_payload_stateElements_1;
    partialRound_tempInput_delay_24_payload_stateElements_2 <= partialRound_tempInput_delay_23_payload_stateElements_2;
    partialRound_tempInput_delay_24_payload_stateElements_3 <= partialRound_tempInput_delay_23_payload_stateElements_3;
    partialRound_tempInput_delay_24_payload_stateElements_4 <= partialRound_tempInput_delay_23_payload_stateElements_4;
    partialRound_tempInput_delay_24_payload_stateElements_5 <= partialRound_tempInput_delay_23_payload_stateElements_5;
    partialRound_tempInput_delay_24_payload_stateElements_6 <= partialRound_tempInput_delay_23_payload_stateElements_6;
    partialRound_tempInput_delay_24_payload_stateElements_7 <= partialRound_tempInput_delay_23_payload_stateElements_7;
    partialRound_tempInput_delay_24_payload_stateElements_8 <= partialRound_tempInput_delay_23_payload_stateElements_8;
    partialRound_tempInput_delay_24_payload_stateElements_9 <= partialRound_tempInput_delay_23_payload_stateElements_9;
    partialRound_tempInput_delay_24_payload_stateElements_10 <= partialRound_tempInput_delay_23_payload_stateElements_10;
    partialRound_tempInput_delay_24_payload_stateElements_11 <= partialRound_tempInput_delay_23_payload_stateElements_11;
    partialRound_tempInput_delay_25_valid <= partialRound_tempInput_delay_24_valid;
    partialRound_tempInput_delay_25_payload_isFull <= partialRound_tempInput_delay_24_payload_isFull;
    partialRound_tempInput_delay_25_payload_fullRound <= partialRound_tempInput_delay_24_payload_fullRound;
    partialRound_tempInput_delay_25_payload_partialRound <= partialRound_tempInput_delay_24_payload_partialRound;
    partialRound_tempInput_delay_25_payload_stateSize <= partialRound_tempInput_delay_24_payload_stateSize;
    partialRound_tempInput_delay_25_payload_stateID <= partialRound_tempInput_delay_24_payload_stateID;
    partialRound_tempInput_delay_25_payload_stateElements_0 <= partialRound_tempInput_delay_24_payload_stateElements_0;
    partialRound_tempInput_delay_25_payload_stateElements_1 <= partialRound_tempInput_delay_24_payload_stateElements_1;
    partialRound_tempInput_delay_25_payload_stateElements_2 <= partialRound_tempInput_delay_24_payload_stateElements_2;
    partialRound_tempInput_delay_25_payload_stateElements_3 <= partialRound_tempInput_delay_24_payload_stateElements_3;
    partialRound_tempInput_delay_25_payload_stateElements_4 <= partialRound_tempInput_delay_24_payload_stateElements_4;
    partialRound_tempInput_delay_25_payload_stateElements_5 <= partialRound_tempInput_delay_24_payload_stateElements_5;
    partialRound_tempInput_delay_25_payload_stateElements_6 <= partialRound_tempInput_delay_24_payload_stateElements_6;
    partialRound_tempInput_delay_25_payload_stateElements_7 <= partialRound_tempInput_delay_24_payload_stateElements_7;
    partialRound_tempInput_delay_25_payload_stateElements_8 <= partialRound_tempInput_delay_24_payload_stateElements_8;
    partialRound_tempInput_delay_25_payload_stateElements_9 <= partialRound_tempInput_delay_24_payload_stateElements_9;
    partialRound_tempInput_delay_25_payload_stateElements_10 <= partialRound_tempInput_delay_24_payload_stateElements_10;
    partialRound_tempInput_delay_25_payload_stateElements_11 <= partialRound_tempInput_delay_24_payload_stateElements_11;
    partialRound_tempInput_delay_26_valid <= partialRound_tempInput_delay_25_valid;
    partialRound_tempInput_delay_26_payload_isFull <= partialRound_tempInput_delay_25_payload_isFull;
    partialRound_tempInput_delay_26_payload_fullRound <= partialRound_tempInput_delay_25_payload_fullRound;
    partialRound_tempInput_delay_26_payload_partialRound <= partialRound_tempInput_delay_25_payload_partialRound;
    partialRound_tempInput_delay_26_payload_stateSize <= partialRound_tempInput_delay_25_payload_stateSize;
    partialRound_tempInput_delay_26_payload_stateID <= partialRound_tempInput_delay_25_payload_stateID;
    partialRound_tempInput_delay_26_payload_stateElements_0 <= partialRound_tempInput_delay_25_payload_stateElements_0;
    partialRound_tempInput_delay_26_payload_stateElements_1 <= partialRound_tempInput_delay_25_payload_stateElements_1;
    partialRound_tempInput_delay_26_payload_stateElements_2 <= partialRound_tempInput_delay_25_payload_stateElements_2;
    partialRound_tempInput_delay_26_payload_stateElements_3 <= partialRound_tempInput_delay_25_payload_stateElements_3;
    partialRound_tempInput_delay_26_payload_stateElements_4 <= partialRound_tempInput_delay_25_payload_stateElements_4;
    partialRound_tempInput_delay_26_payload_stateElements_5 <= partialRound_tempInput_delay_25_payload_stateElements_5;
    partialRound_tempInput_delay_26_payload_stateElements_6 <= partialRound_tempInput_delay_25_payload_stateElements_6;
    partialRound_tempInput_delay_26_payload_stateElements_7 <= partialRound_tempInput_delay_25_payload_stateElements_7;
    partialRound_tempInput_delay_26_payload_stateElements_8 <= partialRound_tempInput_delay_25_payload_stateElements_8;
    partialRound_tempInput_delay_26_payload_stateElements_9 <= partialRound_tempInput_delay_25_payload_stateElements_9;
    partialRound_tempInput_delay_26_payload_stateElements_10 <= partialRound_tempInput_delay_25_payload_stateElements_10;
    partialRound_tempInput_delay_26_payload_stateElements_11 <= partialRound_tempInput_delay_25_payload_stateElements_11;
    partialRound_tempInput_delay_27_valid <= partialRound_tempInput_delay_26_valid;
    partialRound_tempInput_delay_27_payload_isFull <= partialRound_tempInput_delay_26_payload_isFull;
    partialRound_tempInput_delay_27_payload_fullRound <= partialRound_tempInput_delay_26_payload_fullRound;
    partialRound_tempInput_delay_27_payload_partialRound <= partialRound_tempInput_delay_26_payload_partialRound;
    partialRound_tempInput_delay_27_payload_stateSize <= partialRound_tempInput_delay_26_payload_stateSize;
    partialRound_tempInput_delay_27_payload_stateID <= partialRound_tempInput_delay_26_payload_stateID;
    partialRound_tempInput_delay_27_payload_stateElements_0 <= partialRound_tempInput_delay_26_payload_stateElements_0;
    partialRound_tempInput_delay_27_payload_stateElements_1 <= partialRound_tempInput_delay_26_payload_stateElements_1;
    partialRound_tempInput_delay_27_payload_stateElements_2 <= partialRound_tempInput_delay_26_payload_stateElements_2;
    partialRound_tempInput_delay_27_payload_stateElements_3 <= partialRound_tempInput_delay_26_payload_stateElements_3;
    partialRound_tempInput_delay_27_payload_stateElements_4 <= partialRound_tempInput_delay_26_payload_stateElements_4;
    partialRound_tempInput_delay_27_payload_stateElements_5 <= partialRound_tempInput_delay_26_payload_stateElements_5;
    partialRound_tempInput_delay_27_payload_stateElements_6 <= partialRound_tempInput_delay_26_payload_stateElements_6;
    partialRound_tempInput_delay_27_payload_stateElements_7 <= partialRound_tempInput_delay_26_payload_stateElements_7;
    partialRound_tempInput_delay_27_payload_stateElements_8 <= partialRound_tempInput_delay_26_payload_stateElements_8;
    partialRound_tempInput_delay_27_payload_stateElements_9 <= partialRound_tempInput_delay_26_payload_stateElements_9;
    partialRound_tempInput_delay_27_payload_stateElements_10 <= partialRound_tempInput_delay_26_payload_stateElements_10;
    partialRound_tempInput_delay_27_payload_stateElements_11 <= partialRound_tempInput_delay_26_payload_stateElements_11;
    partialRound_tempInput_delay_28_valid <= partialRound_tempInput_delay_27_valid;
    partialRound_tempInput_delay_28_payload_isFull <= partialRound_tempInput_delay_27_payload_isFull;
    partialRound_tempInput_delay_28_payload_fullRound <= partialRound_tempInput_delay_27_payload_fullRound;
    partialRound_tempInput_delay_28_payload_partialRound <= partialRound_tempInput_delay_27_payload_partialRound;
    partialRound_tempInput_delay_28_payload_stateSize <= partialRound_tempInput_delay_27_payload_stateSize;
    partialRound_tempInput_delay_28_payload_stateID <= partialRound_tempInput_delay_27_payload_stateID;
    partialRound_tempInput_delay_28_payload_stateElements_0 <= partialRound_tempInput_delay_27_payload_stateElements_0;
    partialRound_tempInput_delay_28_payload_stateElements_1 <= partialRound_tempInput_delay_27_payload_stateElements_1;
    partialRound_tempInput_delay_28_payload_stateElements_2 <= partialRound_tempInput_delay_27_payload_stateElements_2;
    partialRound_tempInput_delay_28_payload_stateElements_3 <= partialRound_tempInput_delay_27_payload_stateElements_3;
    partialRound_tempInput_delay_28_payload_stateElements_4 <= partialRound_tempInput_delay_27_payload_stateElements_4;
    partialRound_tempInput_delay_28_payload_stateElements_5 <= partialRound_tempInput_delay_27_payload_stateElements_5;
    partialRound_tempInput_delay_28_payload_stateElements_6 <= partialRound_tempInput_delay_27_payload_stateElements_6;
    partialRound_tempInput_delay_28_payload_stateElements_7 <= partialRound_tempInput_delay_27_payload_stateElements_7;
    partialRound_tempInput_delay_28_payload_stateElements_8 <= partialRound_tempInput_delay_27_payload_stateElements_8;
    partialRound_tempInput_delay_28_payload_stateElements_9 <= partialRound_tempInput_delay_27_payload_stateElements_9;
    partialRound_tempInput_delay_28_payload_stateElements_10 <= partialRound_tempInput_delay_27_payload_stateElements_10;
    partialRound_tempInput_delay_28_payload_stateElements_11 <= partialRound_tempInput_delay_27_payload_stateElements_11;
    partialRound_tempInput_delay_29_valid <= partialRound_tempInput_delay_28_valid;
    partialRound_tempInput_delay_29_payload_isFull <= partialRound_tempInput_delay_28_payload_isFull;
    partialRound_tempInput_delay_29_payload_fullRound <= partialRound_tempInput_delay_28_payload_fullRound;
    partialRound_tempInput_delay_29_payload_partialRound <= partialRound_tempInput_delay_28_payload_partialRound;
    partialRound_tempInput_delay_29_payload_stateSize <= partialRound_tempInput_delay_28_payload_stateSize;
    partialRound_tempInput_delay_29_payload_stateID <= partialRound_tempInput_delay_28_payload_stateID;
    partialRound_tempInput_delay_29_payload_stateElements_0 <= partialRound_tempInput_delay_28_payload_stateElements_0;
    partialRound_tempInput_delay_29_payload_stateElements_1 <= partialRound_tempInput_delay_28_payload_stateElements_1;
    partialRound_tempInput_delay_29_payload_stateElements_2 <= partialRound_tempInput_delay_28_payload_stateElements_2;
    partialRound_tempInput_delay_29_payload_stateElements_3 <= partialRound_tempInput_delay_28_payload_stateElements_3;
    partialRound_tempInput_delay_29_payload_stateElements_4 <= partialRound_tempInput_delay_28_payload_stateElements_4;
    partialRound_tempInput_delay_29_payload_stateElements_5 <= partialRound_tempInput_delay_28_payload_stateElements_5;
    partialRound_tempInput_delay_29_payload_stateElements_6 <= partialRound_tempInput_delay_28_payload_stateElements_6;
    partialRound_tempInput_delay_29_payload_stateElements_7 <= partialRound_tempInput_delay_28_payload_stateElements_7;
    partialRound_tempInput_delay_29_payload_stateElements_8 <= partialRound_tempInput_delay_28_payload_stateElements_8;
    partialRound_tempInput_delay_29_payload_stateElements_9 <= partialRound_tempInput_delay_28_payload_stateElements_9;
    partialRound_tempInput_delay_29_payload_stateElements_10 <= partialRound_tempInput_delay_28_payload_stateElements_10;
    partialRound_tempInput_delay_29_payload_stateElements_11 <= partialRound_tempInput_delay_28_payload_stateElements_11;
    partialRound_tempInput_delay_30_valid <= partialRound_tempInput_delay_29_valid;
    partialRound_tempInput_delay_30_payload_isFull <= partialRound_tempInput_delay_29_payload_isFull;
    partialRound_tempInput_delay_30_payload_fullRound <= partialRound_tempInput_delay_29_payload_fullRound;
    partialRound_tempInput_delay_30_payload_partialRound <= partialRound_tempInput_delay_29_payload_partialRound;
    partialRound_tempInput_delay_30_payload_stateSize <= partialRound_tempInput_delay_29_payload_stateSize;
    partialRound_tempInput_delay_30_payload_stateID <= partialRound_tempInput_delay_29_payload_stateID;
    partialRound_tempInput_delay_30_payload_stateElements_0 <= partialRound_tempInput_delay_29_payload_stateElements_0;
    partialRound_tempInput_delay_30_payload_stateElements_1 <= partialRound_tempInput_delay_29_payload_stateElements_1;
    partialRound_tempInput_delay_30_payload_stateElements_2 <= partialRound_tempInput_delay_29_payload_stateElements_2;
    partialRound_tempInput_delay_30_payload_stateElements_3 <= partialRound_tempInput_delay_29_payload_stateElements_3;
    partialRound_tempInput_delay_30_payload_stateElements_4 <= partialRound_tempInput_delay_29_payload_stateElements_4;
    partialRound_tempInput_delay_30_payload_stateElements_5 <= partialRound_tempInput_delay_29_payload_stateElements_5;
    partialRound_tempInput_delay_30_payload_stateElements_6 <= partialRound_tempInput_delay_29_payload_stateElements_6;
    partialRound_tempInput_delay_30_payload_stateElements_7 <= partialRound_tempInput_delay_29_payload_stateElements_7;
    partialRound_tempInput_delay_30_payload_stateElements_8 <= partialRound_tempInput_delay_29_payload_stateElements_8;
    partialRound_tempInput_delay_30_payload_stateElements_9 <= partialRound_tempInput_delay_29_payload_stateElements_9;
    partialRound_tempInput_delay_30_payload_stateElements_10 <= partialRound_tempInput_delay_29_payload_stateElements_10;
    partialRound_tempInput_delay_30_payload_stateElements_11 <= partialRound_tempInput_delay_29_payload_stateElements_11;
    partialRound_tempInput_delay_31_valid <= partialRound_tempInput_delay_30_valid;
    partialRound_tempInput_delay_31_payload_isFull <= partialRound_tempInput_delay_30_payload_isFull;
    partialRound_tempInput_delay_31_payload_fullRound <= partialRound_tempInput_delay_30_payload_fullRound;
    partialRound_tempInput_delay_31_payload_partialRound <= partialRound_tempInput_delay_30_payload_partialRound;
    partialRound_tempInput_delay_31_payload_stateSize <= partialRound_tempInput_delay_30_payload_stateSize;
    partialRound_tempInput_delay_31_payload_stateID <= partialRound_tempInput_delay_30_payload_stateID;
    partialRound_tempInput_delay_31_payload_stateElements_0 <= partialRound_tempInput_delay_30_payload_stateElements_0;
    partialRound_tempInput_delay_31_payload_stateElements_1 <= partialRound_tempInput_delay_30_payload_stateElements_1;
    partialRound_tempInput_delay_31_payload_stateElements_2 <= partialRound_tempInput_delay_30_payload_stateElements_2;
    partialRound_tempInput_delay_31_payload_stateElements_3 <= partialRound_tempInput_delay_30_payload_stateElements_3;
    partialRound_tempInput_delay_31_payload_stateElements_4 <= partialRound_tempInput_delay_30_payload_stateElements_4;
    partialRound_tempInput_delay_31_payload_stateElements_5 <= partialRound_tempInput_delay_30_payload_stateElements_5;
    partialRound_tempInput_delay_31_payload_stateElements_6 <= partialRound_tempInput_delay_30_payload_stateElements_6;
    partialRound_tempInput_delay_31_payload_stateElements_7 <= partialRound_tempInput_delay_30_payload_stateElements_7;
    partialRound_tempInput_delay_31_payload_stateElements_8 <= partialRound_tempInput_delay_30_payload_stateElements_8;
    partialRound_tempInput_delay_31_payload_stateElements_9 <= partialRound_tempInput_delay_30_payload_stateElements_9;
    partialRound_tempInput_delay_31_payload_stateElements_10 <= partialRound_tempInput_delay_30_payload_stateElements_10;
    partialRound_tempInput_delay_31_payload_stateElements_11 <= partialRound_tempInput_delay_30_payload_stateElements_11;
    partialRound_tempInput_delay_32_valid <= partialRound_tempInput_delay_31_valid;
    partialRound_tempInput_delay_32_payload_isFull <= partialRound_tempInput_delay_31_payload_isFull;
    partialRound_tempInput_delay_32_payload_fullRound <= partialRound_tempInput_delay_31_payload_fullRound;
    partialRound_tempInput_delay_32_payload_partialRound <= partialRound_tempInput_delay_31_payload_partialRound;
    partialRound_tempInput_delay_32_payload_stateSize <= partialRound_tempInput_delay_31_payload_stateSize;
    partialRound_tempInput_delay_32_payload_stateID <= partialRound_tempInput_delay_31_payload_stateID;
    partialRound_tempInput_delay_32_payload_stateElements_0 <= partialRound_tempInput_delay_31_payload_stateElements_0;
    partialRound_tempInput_delay_32_payload_stateElements_1 <= partialRound_tempInput_delay_31_payload_stateElements_1;
    partialRound_tempInput_delay_32_payload_stateElements_2 <= partialRound_tempInput_delay_31_payload_stateElements_2;
    partialRound_tempInput_delay_32_payload_stateElements_3 <= partialRound_tempInput_delay_31_payload_stateElements_3;
    partialRound_tempInput_delay_32_payload_stateElements_4 <= partialRound_tempInput_delay_31_payload_stateElements_4;
    partialRound_tempInput_delay_32_payload_stateElements_5 <= partialRound_tempInput_delay_31_payload_stateElements_5;
    partialRound_tempInput_delay_32_payload_stateElements_6 <= partialRound_tempInput_delay_31_payload_stateElements_6;
    partialRound_tempInput_delay_32_payload_stateElements_7 <= partialRound_tempInput_delay_31_payload_stateElements_7;
    partialRound_tempInput_delay_32_payload_stateElements_8 <= partialRound_tempInput_delay_31_payload_stateElements_8;
    partialRound_tempInput_delay_32_payload_stateElements_9 <= partialRound_tempInput_delay_31_payload_stateElements_9;
    partialRound_tempInput_delay_32_payload_stateElements_10 <= partialRound_tempInput_delay_31_payload_stateElements_10;
    partialRound_tempInput_delay_32_payload_stateElements_11 <= partialRound_tempInput_delay_31_payload_stateElements_11;
    partialRound_tempInput_delay_33_valid <= partialRound_tempInput_delay_32_valid;
    partialRound_tempInput_delay_33_payload_isFull <= partialRound_tempInput_delay_32_payload_isFull;
    partialRound_tempInput_delay_33_payload_fullRound <= partialRound_tempInput_delay_32_payload_fullRound;
    partialRound_tempInput_delay_33_payload_partialRound <= partialRound_tempInput_delay_32_payload_partialRound;
    partialRound_tempInput_delay_33_payload_stateSize <= partialRound_tempInput_delay_32_payload_stateSize;
    partialRound_tempInput_delay_33_payload_stateID <= partialRound_tempInput_delay_32_payload_stateID;
    partialRound_tempInput_delay_33_payload_stateElements_0 <= partialRound_tempInput_delay_32_payload_stateElements_0;
    partialRound_tempInput_delay_33_payload_stateElements_1 <= partialRound_tempInput_delay_32_payload_stateElements_1;
    partialRound_tempInput_delay_33_payload_stateElements_2 <= partialRound_tempInput_delay_32_payload_stateElements_2;
    partialRound_tempInput_delay_33_payload_stateElements_3 <= partialRound_tempInput_delay_32_payload_stateElements_3;
    partialRound_tempInput_delay_33_payload_stateElements_4 <= partialRound_tempInput_delay_32_payload_stateElements_4;
    partialRound_tempInput_delay_33_payload_stateElements_5 <= partialRound_tempInput_delay_32_payload_stateElements_5;
    partialRound_tempInput_delay_33_payload_stateElements_6 <= partialRound_tempInput_delay_32_payload_stateElements_6;
    partialRound_tempInput_delay_33_payload_stateElements_7 <= partialRound_tempInput_delay_32_payload_stateElements_7;
    partialRound_tempInput_delay_33_payload_stateElements_8 <= partialRound_tempInput_delay_32_payload_stateElements_8;
    partialRound_tempInput_delay_33_payload_stateElements_9 <= partialRound_tempInput_delay_32_payload_stateElements_9;
    partialRound_tempInput_delay_33_payload_stateElements_10 <= partialRound_tempInput_delay_32_payload_stateElements_10;
    partialRound_tempInput_delay_33_payload_stateElements_11 <= partialRound_tempInput_delay_32_payload_stateElements_11;
    partialRound_tempInput_delay_34_valid <= partialRound_tempInput_delay_33_valid;
    partialRound_tempInput_delay_34_payload_isFull <= partialRound_tempInput_delay_33_payload_isFull;
    partialRound_tempInput_delay_34_payload_fullRound <= partialRound_tempInput_delay_33_payload_fullRound;
    partialRound_tempInput_delay_34_payload_partialRound <= partialRound_tempInput_delay_33_payload_partialRound;
    partialRound_tempInput_delay_34_payload_stateSize <= partialRound_tempInput_delay_33_payload_stateSize;
    partialRound_tempInput_delay_34_payload_stateID <= partialRound_tempInput_delay_33_payload_stateID;
    partialRound_tempInput_delay_34_payload_stateElements_0 <= partialRound_tempInput_delay_33_payload_stateElements_0;
    partialRound_tempInput_delay_34_payload_stateElements_1 <= partialRound_tempInput_delay_33_payload_stateElements_1;
    partialRound_tempInput_delay_34_payload_stateElements_2 <= partialRound_tempInput_delay_33_payload_stateElements_2;
    partialRound_tempInput_delay_34_payload_stateElements_3 <= partialRound_tempInput_delay_33_payload_stateElements_3;
    partialRound_tempInput_delay_34_payload_stateElements_4 <= partialRound_tempInput_delay_33_payload_stateElements_4;
    partialRound_tempInput_delay_34_payload_stateElements_5 <= partialRound_tempInput_delay_33_payload_stateElements_5;
    partialRound_tempInput_delay_34_payload_stateElements_6 <= partialRound_tempInput_delay_33_payload_stateElements_6;
    partialRound_tempInput_delay_34_payload_stateElements_7 <= partialRound_tempInput_delay_33_payload_stateElements_7;
    partialRound_tempInput_delay_34_payload_stateElements_8 <= partialRound_tempInput_delay_33_payload_stateElements_8;
    partialRound_tempInput_delay_34_payload_stateElements_9 <= partialRound_tempInput_delay_33_payload_stateElements_9;
    partialRound_tempInput_delay_34_payload_stateElements_10 <= partialRound_tempInput_delay_33_payload_stateElements_10;
    partialRound_tempInput_delay_34_payload_stateElements_11 <= partialRound_tempInput_delay_33_payload_stateElements_11;
    partialRound_tempInput_delay_35_valid <= partialRound_tempInput_delay_34_valid;
    partialRound_tempInput_delay_35_payload_isFull <= partialRound_tempInput_delay_34_payload_isFull;
    partialRound_tempInput_delay_35_payload_fullRound <= partialRound_tempInput_delay_34_payload_fullRound;
    partialRound_tempInput_delay_35_payload_partialRound <= partialRound_tempInput_delay_34_payload_partialRound;
    partialRound_tempInput_delay_35_payload_stateSize <= partialRound_tempInput_delay_34_payload_stateSize;
    partialRound_tempInput_delay_35_payload_stateID <= partialRound_tempInput_delay_34_payload_stateID;
    partialRound_tempInput_delay_35_payload_stateElements_0 <= partialRound_tempInput_delay_34_payload_stateElements_0;
    partialRound_tempInput_delay_35_payload_stateElements_1 <= partialRound_tempInput_delay_34_payload_stateElements_1;
    partialRound_tempInput_delay_35_payload_stateElements_2 <= partialRound_tempInput_delay_34_payload_stateElements_2;
    partialRound_tempInput_delay_35_payload_stateElements_3 <= partialRound_tempInput_delay_34_payload_stateElements_3;
    partialRound_tempInput_delay_35_payload_stateElements_4 <= partialRound_tempInput_delay_34_payload_stateElements_4;
    partialRound_tempInput_delay_35_payload_stateElements_5 <= partialRound_tempInput_delay_34_payload_stateElements_5;
    partialRound_tempInput_delay_35_payload_stateElements_6 <= partialRound_tempInput_delay_34_payload_stateElements_6;
    partialRound_tempInput_delay_35_payload_stateElements_7 <= partialRound_tempInput_delay_34_payload_stateElements_7;
    partialRound_tempInput_delay_35_payload_stateElements_8 <= partialRound_tempInput_delay_34_payload_stateElements_8;
    partialRound_tempInput_delay_35_payload_stateElements_9 <= partialRound_tempInput_delay_34_payload_stateElements_9;
    partialRound_tempInput_delay_35_payload_stateElements_10 <= partialRound_tempInput_delay_34_payload_stateElements_10;
    partialRound_tempInput_delay_35_payload_stateElements_11 <= partialRound_tempInput_delay_34_payload_stateElements_11;
    partialRound_tempInput_delay_36_valid <= partialRound_tempInput_delay_35_valid;
    partialRound_tempInput_delay_36_payload_isFull <= partialRound_tempInput_delay_35_payload_isFull;
    partialRound_tempInput_delay_36_payload_fullRound <= partialRound_tempInput_delay_35_payload_fullRound;
    partialRound_tempInput_delay_36_payload_partialRound <= partialRound_tempInput_delay_35_payload_partialRound;
    partialRound_tempInput_delay_36_payload_stateSize <= partialRound_tempInput_delay_35_payload_stateSize;
    partialRound_tempInput_delay_36_payload_stateID <= partialRound_tempInput_delay_35_payload_stateID;
    partialRound_tempInput_delay_36_payload_stateElements_0 <= partialRound_tempInput_delay_35_payload_stateElements_0;
    partialRound_tempInput_delay_36_payload_stateElements_1 <= partialRound_tempInput_delay_35_payload_stateElements_1;
    partialRound_tempInput_delay_36_payload_stateElements_2 <= partialRound_tempInput_delay_35_payload_stateElements_2;
    partialRound_tempInput_delay_36_payload_stateElements_3 <= partialRound_tempInput_delay_35_payload_stateElements_3;
    partialRound_tempInput_delay_36_payload_stateElements_4 <= partialRound_tempInput_delay_35_payload_stateElements_4;
    partialRound_tempInput_delay_36_payload_stateElements_5 <= partialRound_tempInput_delay_35_payload_stateElements_5;
    partialRound_tempInput_delay_36_payload_stateElements_6 <= partialRound_tempInput_delay_35_payload_stateElements_6;
    partialRound_tempInput_delay_36_payload_stateElements_7 <= partialRound_tempInput_delay_35_payload_stateElements_7;
    partialRound_tempInput_delay_36_payload_stateElements_8 <= partialRound_tempInput_delay_35_payload_stateElements_8;
    partialRound_tempInput_delay_36_payload_stateElements_9 <= partialRound_tempInput_delay_35_payload_stateElements_9;
    partialRound_tempInput_delay_36_payload_stateElements_10 <= partialRound_tempInput_delay_35_payload_stateElements_10;
    partialRound_tempInput_delay_36_payload_stateElements_11 <= partialRound_tempInput_delay_35_payload_stateElements_11;
    partialRound_tempInput_delay_37_valid <= partialRound_tempInput_delay_36_valid;
    partialRound_tempInput_delay_37_payload_isFull <= partialRound_tempInput_delay_36_payload_isFull;
    partialRound_tempInput_delay_37_payload_fullRound <= partialRound_tempInput_delay_36_payload_fullRound;
    partialRound_tempInput_delay_37_payload_partialRound <= partialRound_tempInput_delay_36_payload_partialRound;
    partialRound_tempInput_delay_37_payload_stateSize <= partialRound_tempInput_delay_36_payload_stateSize;
    partialRound_tempInput_delay_37_payload_stateID <= partialRound_tempInput_delay_36_payload_stateID;
    partialRound_tempInput_delay_37_payload_stateElements_0 <= partialRound_tempInput_delay_36_payload_stateElements_0;
    partialRound_tempInput_delay_37_payload_stateElements_1 <= partialRound_tempInput_delay_36_payload_stateElements_1;
    partialRound_tempInput_delay_37_payload_stateElements_2 <= partialRound_tempInput_delay_36_payload_stateElements_2;
    partialRound_tempInput_delay_37_payload_stateElements_3 <= partialRound_tempInput_delay_36_payload_stateElements_3;
    partialRound_tempInput_delay_37_payload_stateElements_4 <= partialRound_tempInput_delay_36_payload_stateElements_4;
    partialRound_tempInput_delay_37_payload_stateElements_5 <= partialRound_tempInput_delay_36_payload_stateElements_5;
    partialRound_tempInput_delay_37_payload_stateElements_6 <= partialRound_tempInput_delay_36_payload_stateElements_6;
    partialRound_tempInput_delay_37_payload_stateElements_7 <= partialRound_tempInput_delay_36_payload_stateElements_7;
    partialRound_tempInput_delay_37_payload_stateElements_8 <= partialRound_tempInput_delay_36_payload_stateElements_8;
    partialRound_tempInput_delay_37_payload_stateElements_9 <= partialRound_tempInput_delay_36_payload_stateElements_9;
    partialRound_tempInput_delay_37_payload_stateElements_10 <= partialRound_tempInput_delay_36_payload_stateElements_10;
    partialRound_tempInput_delay_37_payload_stateElements_11 <= partialRound_tempInput_delay_36_payload_stateElements_11;
    partialRound_tempInput_delay_38_valid <= partialRound_tempInput_delay_37_valid;
    partialRound_tempInput_delay_38_payload_isFull <= partialRound_tempInput_delay_37_payload_isFull;
    partialRound_tempInput_delay_38_payload_fullRound <= partialRound_tempInput_delay_37_payload_fullRound;
    partialRound_tempInput_delay_38_payload_partialRound <= partialRound_tempInput_delay_37_payload_partialRound;
    partialRound_tempInput_delay_38_payload_stateSize <= partialRound_tempInput_delay_37_payload_stateSize;
    partialRound_tempInput_delay_38_payload_stateID <= partialRound_tempInput_delay_37_payload_stateID;
    partialRound_tempInput_delay_38_payload_stateElements_0 <= partialRound_tempInput_delay_37_payload_stateElements_0;
    partialRound_tempInput_delay_38_payload_stateElements_1 <= partialRound_tempInput_delay_37_payload_stateElements_1;
    partialRound_tempInput_delay_38_payload_stateElements_2 <= partialRound_tempInput_delay_37_payload_stateElements_2;
    partialRound_tempInput_delay_38_payload_stateElements_3 <= partialRound_tempInput_delay_37_payload_stateElements_3;
    partialRound_tempInput_delay_38_payload_stateElements_4 <= partialRound_tempInput_delay_37_payload_stateElements_4;
    partialRound_tempInput_delay_38_payload_stateElements_5 <= partialRound_tempInput_delay_37_payload_stateElements_5;
    partialRound_tempInput_delay_38_payload_stateElements_6 <= partialRound_tempInput_delay_37_payload_stateElements_6;
    partialRound_tempInput_delay_38_payload_stateElements_7 <= partialRound_tempInput_delay_37_payload_stateElements_7;
    partialRound_tempInput_delay_38_payload_stateElements_8 <= partialRound_tempInput_delay_37_payload_stateElements_8;
    partialRound_tempInput_delay_38_payload_stateElements_9 <= partialRound_tempInput_delay_37_payload_stateElements_9;
    partialRound_tempInput_delay_38_payload_stateElements_10 <= partialRound_tempInput_delay_37_payload_stateElements_10;
    partialRound_tempInput_delay_38_payload_stateElements_11 <= partialRound_tempInput_delay_37_payload_stateElements_11;
    partialRound_tempInput_delay_39_valid <= partialRound_tempInput_delay_38_valid;
    partialRound_tempInput_delay_39_payload_isFull <= partialRound_tempInput_delay_38_payload_isFull;
    partialRound_tempInput_delay_39_payload_fullRound <= partialRound_tempInput_delay_38_payload_fullRound;
    partialRound_tempInput_delay_39_payload_partialRound <= partialRound_tempInput_delay_38_payload_partialRound;
    partialRound_tempInput_delay_39_payload_stateSize <= partialRound_tempInput_delay_38_payload_stateSize;
    partialRound_tempInput_delay_39_payload_stateID <= partialRound_tempInput_delay_38_payload_stateID;
    partialRound_tempInput_delay_39_payload_stateElements_0 <= partialRound_tempInput_delay_38_payload_stateElements_0;
    partialRound_tempInput_delay_39_payload_stateElements_1 <= partialRound_tempInput_delay_38_payload_stateElements_1;
    partialRound_tempInput_delay_39_payload_stateElements_2 <= partialRound_tempInput_delay_38_payload_stateElements_2;
    partialRound_tempInput_delay_39_payload_stateElements_3 <= partialRound_tempInput_delay_38_payload_stateElements_3;
    partialRound_tempInput_delay_39_payload_stateElements_4 <= partialRound_tempInput_delay_38_payload_stateElements_4;
    partialRound_tempInput_delay_39_payload_stateElements_5 <= partialRound_tempInput_delay_38_payload_stateElements_5;
    partialRound_tempInput_delay_39_payload_stateElements_6 <= partialRound_tempInput_delay_38_payload_stateElements_6;
    partialRound_tempInput_delay_39_payload_stateElements_7 <= partialRound_tempInput_delay_38_payload_stateElements_7;
    partialRound_tempInput_delay_39_payload_stateElements_8 <= partialRound_tempInput_delay_38_payload_stateElements_8;
    partialRound_tempInput_delay_39_payload_stateElements_9 <= partialRound_tempInput_delay_38_payload_stateElements_9;
    partialRound_tempInput_delay_39_payload_stateElements_10 <= partialRound_tempInput_delay_38_payload_stateElements_10;
    partialRound_tempInput_delay_39_payload_stateElements_11 <= partialRound_tempInput_delay_38_payload_stateElements_11;
    partialRound_tempInput_delay_40_valid <= partialRound_tempInput_delay_39_valid;
    partialRound_tempInput_delay_40_payload_isFull <= partialRound_tempInput_delay_39_payload_isFull;
    partialRound_tempInput_delay_40_payload_fullRound <= partialRound_tempInput_delay_39_payload_fullRound;
    partialRound_tempInput_delay_40_payload_partialRound <= partialRound_tempInput_delay_39_payload_partialRound;
    partialRound_tempInput_delay_40_payload_stateSize <= partialRound_tempInput_delay_39_payload_stateSize;
    partialRound_tempInput_delay_40_payload_stateID <= partialRound_tempInput_delay_39_payload_stateID;
    partialRound_tempInput_delay_40_payload_stateElements_0 <= partialRound_tempInput_delay_39_payload_stateElements_0;
    partialRound_tempInput_delay_40_payload_stateElements_1 <= partialRound_tempInput_delay_39_payload_stateElements_1;
    partialRound_tempInput_delay_40_payload_stateElements_2 <= partialRound_tempInput_delay_39_payload_stateElements_2;
    partialRound_tempInput_delay_40_payload_stateElements_3 <= partialRound_tempInput_delay_39_payload_stateElements_3;
    partialRound_tempInput_delay_40_payload_stateElements_4 <= partialRound_tempInput_delay_39_payload_stateElements_4;
    partialRound_tempInput_delay_40_payload_stateElements_5 <= partialRound_tempInput_delay_39_payload_stateElements_5;
    partialRound_tempInput_delay_40_payload_stateElements_6 <= partialRound_tempInput_delay_39_payload_stateElements_6;
    partialRound_tempInput_delay_40_payload_stateElements_7 <= partialRound_tempInput_delay_39_payload_stateElements_7;
    partialRound_tempInput_delay_40_payload_stateElements_8 <= partialRound_tempInput_delay_39_payload_stateElements_8;
    partialRound_tempInput_delay_40_payload_stateElements_9 <= partialRound_tempInput_delay_39_payload_stateElements_9;
    partialRound_tempInput_delay_40_payload_stateElements_10 <= partialRound_tempInput_delay_39_payload_stateElements_10;
    partialRound_tempInput_delay_40_payload_stateElements_11 <= partialRound_tempInput_delay_39_payload_stateElements_11;
    partialRound_tempInput_delay_41_valid <= partialRound_tempInput_delay_40_valid;
    partialRound_tempInput_delay_41_payload_isFull <= partialRound_tempInput_delay_40_payload_isFull;
    partialRound_tempInput_delay_41_payload_fullRound <= partialRound_tempInput_delay_40_payload_fullRound;
    partialRound_tempInput_delay_41_payload_partialRound <= partialRound_tempInput_delay_40_payload_partialRound;
    partialRound_tempInput_delay_41_payload_stateSize <= partialRound_tempInput_delay_40_payload_stateSize;
    partialRound_tempInput_delay_41_payload_stateID <= partialRound_tempInput_delay_40_payload_stateID;
    partialRound_tempInput_delay_41_payload_stateElements_0 <= partialRound_tempInput_delay_40_payload_stateElements_0;
    partialRound_tempInput_delay_41_payload_stateElements_1 <= partialRound_tempInput_delay_40_payload_stateElements_1;
    partialRound_tempInput_delay_41_payload_stateElements_2 <= partialRound_tempInput_delay_40_payload_stateElements_2;
    partialRound_tempInput_delay_41_payload_stateElements_3 <= partialRound_tempInput_delay_40_payload_stateElements_3;
    partialRound_tempInput_delay_41_payload_stateElements_4 <= partialRound_tempInput_delay_40_payload_stateElements_4;
    partialRound_tempInput_delay_41_payload_stateElements_5 <= partialRound_tempInput_delay_40_payload_stateElements_5;
    partialRound_tempInput_delay_41_payload_stateElements_6 <= partialRound_tempInput_delay_40_payload_stateElements_6;
    partialRound_tempInput_delay_41_payload_stateElements_7 <= partialRound_tempInput_delay_40_payload_stateElements_7;
    partialRound_tempInput_delay_41_payload_stateElements_8 <= partialRound_tempInput_delay_40_payload_stateElements_8;
    partialRound_tempInput_delay_41_payload_stateElements_9 <= partialRound_tempInput_delay_40_payload_stateElements_9;
    partialRound_tempInput_delay_41_payload_stateElements_10 <= partialRound_tempInput_delay_40_payload_stateElements_10;
    partialRound_tempInput_delay_41_payload_stateElements_11 <= partialRound_tempInput_delay_40_payload_stateElements_11;
    partialRound_tempInput_delay_42_valid <= partialRound_tempInput_delay_41_valid;
    partialRound_tempInput_delay_42_payload_isFull <= partialRound_tempInput_delay_41_payload_isFull;
    partialRound_tempInput_delay_42_payload_fullRound <= partialRound_tempInput_delay_41_payload_fullRound;
    partialRound_tempInput_delay_42_payload_partialRound <= partialRound_tempInput_delay_41_payload_partialRound;
    partialRound_tempInput_delay_42_payload_stateSize <= partialRound_tempInput_delay_41_payload_stateSize;
    partialRound_tempInput_delay_42_payload_stateID <= partialRound_tempInput_delay_41_payload_stateID;
    partialRound_tempInput_delay_42_payload_stateElements_0 <= partialRound_tempInput_delay_41_payload_stateElements_0;
    partialRound_tempInput_delay_42_payload_stateElements_1 <= partialRound_tempInput_delay_41_payload_stateElements_1;
    partialRound_tempInput_delay_42_payload_stateElements_2 <= partialRound_tempInput_delay_41_payload_stateElements_2;
    partialRound_tempInput_delay_42_payload_stateElements_3 <= partialRound_tempInput_delay_41_payload_stateElements_3;
    partialRound_tempInput_delay_42_payload_stateElements_4 <= partialRound_tempInput_delay_41_payload_stateElements_4;
    partialRound_tempInput_delay_42_payload_stateElements_5 <= partialRound_tempInput_delay_41_payload_stateElements_5;
    partialRound_tempInput_delay_42_payload_stateElements_6 <= partialRound_tempInput_delay_41_payload_stateElements_6;
    partialRound_tempInput_delay_42_payload_stateElements_7 <= partialRound_tempInput_delay_41_payload_stateElements_7;
    partialRound_tempInput_delay_42_payload_stateElements_8 <= partialRound_tempInput_delay_41_payload_stateElements_8;
    partialRound_tempInput_delay_42_payload_stateElements_9 <= partialRound_tempInput_delay_41_payload_stateElements_9;
    partialRound_tempInput_delay_42_payload_stateElements_10 <= partialRound_tempInput_delay_41_payload_stateElements_10;
    partialRound_tempInput_delay_42_payload_stateElements_11 <= partialRound_tempInput_delay_41_payload_stateElements_11;
    partialRound_tempInput_delay_43_valid <= partialRound_tempInput_delay_42_valid;
    partialRound_tempInput_delay_43_payload_isFull <= partialRound_tempInput_delay_42_payload_isFull;
    partialRound_tempInput_delay_43_payload_fullRound <= partialRound_tempInput_delay_42_payload_fullRound;
    partialRound_tempInput_delay_43_payload_partialRound <= partialRound_tempInput_delay_42_payload_partialRound;
    partialRound_tempInput_delay_43_payload_stateSize <= partialRound_tempInput_delay_42_payload_stateSize;
    partialRound_tempInput_delay_43_payload_stateID <= partialRound_tempInput_delay_42_payload_stateID;
    partialRound_tempInput_delay_43_payload_stateElements_0 <= partialRound_tempInput_delay_42_payload_stateElements_0;
    partialRound_tempInput_delay_43_payload_stateElements_1 <= partialRound_tempInput_delay_42_payload_stateElements_1;
    partialRound_tempInput_delay_43_payload_stateElements_2 <= partialRound_tempInput_delay_42_payload_stateElements_2;
    partialRound_tempInput_delay_43_payload_stateElements_3 <= partialRound_tempInput_delay_42_payload_stateElements_3;
    partialRound_tempInput_delay_43_payload_stateElements_4 <= partialRound_tempInput_delay_42_payload_stateElements_4;
    partialRound_tempInput_delay_43_payload_stateElements_5 <= partialRound_tempInput_delay_42_payload_stateElements_5;
    partialRound_tempInput_delay_43_payload_stateElements_6 <= partialRound_tempInput_delay_42_payload_stateElements_6;
    partialRound_tempInput_delay_43_payload_stateElements_7 <= partialRound_tempInput_delay_42_payload_stateElements_7;
    partialRound_tempInput_delay_43_payload_stateElements_8 <= partialRound_tempInput_delay_42_payload_stateElements_8;
    partialRound_tempInput_delay_43_payload_stateElements_9 <= partialRound_tempInput_delay_42_payload_stateElements_9;
    partialRound_tempInput_delay_43_payload_stateElements_10 <= partialRound_tempInput_delay_42_payload_stateElements_10;
    partialRound_tempInput_delay_43_payload_stateElements_11 <= partialRound_tempInput_delay_42_payload_stateElements_11;
    partialRound_tempInput_delay_44_valid <= partialRound_tempInput_delay_43_valid;
    partialRound_tempInput_delay_44_payload_isFull <= partialRound_tempInput_delay_43_payload_isFull;
    partialRound_tempInput_delay_44_payload_fullRound <= partialRound_tempInput_delay_43_payload_fullRound;
    partialRound_tempInput_delay_44_payload_partialRound <= partialRound_tempInput_delay_43_payload_partialRound;
    partialRound_tempInput_delay_44_payload_stateSize <= partialRound_tempInput_delay_43_payload_stateSize;
    partialRound_tempInput_delay_44_payload_stateID <= partialRound_tempInput_delay_43_payload_stateID;
    partialRound_tempInput_delay_44_payload_stateElements_0 <= partialRound_tempInput_delay_43_payload_stateElements_0;
    partialRound_tempInput_delay_44_payload_stateElements_1 <= partialRound_tempInput_delay_43_payload_stateElements_1;
    partialRound_tempInput_delay_44_payload_stateElements_2 <= partialRound_tempInput_delay_43_payload_stateElements_2;
    partialRound_tempInput_delay_44_payload_stateElements_3 <= partialRound_tempInput_delay_43_payload_stateElements_3;
    partialRound_tempInput_delay_44_payload_stateElements_4 <= partialRound_tempInput_delay_43_payload_stateElements_4;
    partialRound_tempInput_delay_44_payload_stateElements_5 <= partialRound_tempInput_delay_43_payload_stateElements_5;
    partialRound_tempInput_delay_44_payload_stateElements_6 <= partialRound_tempInput_delay_43_payload_stateElements_6;
    partialRound_tempInput_delay_44_payload_stateElements_7 <= partialRound_tempInput_delay_43_payload_stateElements_7;
    partialRound_tempInput_delay_44_payload_stateElements_8 <= partialRound_tempInput_delay_43_payload_stateElements_8;
    partialRound_tempInput_delay_44_payload_stateElements_9 <= partialRound_tempInput_delay_43_payload_stateElements_9;
    partialRound_tempInput_delay_44_payload_stateElements_10 <= partialRound_tempInput_delay_43_payload_stateElements_10;
    partialRound_tempInput_delay_44_payload_stateElements_11 <= partialRound_tempInput_delay_43_payload_stateElements_11;
    partialRound_tempInput_delay_45_valid <= partialRound_tempInput_delay_44_valid;
    partialRound_tempInput_delay_45_payload_isFull <= partialRound_tempInput_delay_44_payload_isFull;
    partialRound_tempInput_delay_45_payload_fullRound <= partialRound_tempInput_delay_44_payload_fullRound;
    partialRound_tempInput_delay_45_payload_partialRound <= partialRound_tempInput_delay_44_payload_partialRound;
    partialRound_tempInput_delay_45_payload_stateSize <= partialRound_tempInput_delay_44_payload_stateSize;
    partialRound_tempInput_delay_45_payload_stateID <= partialRound_tempInput_delay_44_payload_stateID;
    partialRound_tempInput_delay_45_payload_stateElements_0 <= partialRound_tempInput_delay_44_payload_stateElements_0;
    partialRound_tempInput_delay_45_payload_stateElements_1 <= partialRound_tempInput_delay_44_payload_stateElements_1;
    partialRound_tempInput_delay_45_payload_stateElements_2 <= partialRound_tempInput_delay_44_payload_stateElements_2;
    partialRound_tempInput_delay_45_payload_stateElements_3 <= partialRound_tempInput_delay_44_payload_stateElements_3;
    partialRound_tempInput_delay_45_payload_stateElements_4 <= partialRound_tempInput_delay_44_payload_stateElements_4;
    partialRound_tempInput_delay_45_payload_stateElements_5 <= partialRound_tempInput_delay_44_payload_stateElements_5;
    partialRound_tempInput_delay_45_payload_stateElements_6 <= partialRound_tempInput_delay_44_payload_stateElements_6;
    partialRound_tempInput_delay_45_payload_stateElements_7 <= partialRound_tempInput_delay_44_payload_stateElements_7;
    partialRound_tempInput_delay_45_payload_stateElements_8 <= partialRound_tempInput_delay_44_payload_stateElements_8;
    partialRound_tempInput_delay_45_payload_stateElements_9 <= partialRound_tempInput_delay_44_payload_stateElements_9;
    partialRound_tempInput_delay_45_payload_stateElements_10 <= partialRound_tempInput_delay_44_payload_stateElements_10;
    partialRound_tempInput_delay_45_payload_stateElements_11 <= partialRound_tempInput_delay_44_payload_stateElements_11;
    partialRound_tempInput_delay_46_valid <= partialRound_tempInput_delay_45_valid;
    partialRound_tempInput_delay_46_payload_isFull <= partialRound_tempInput_delay_45_payload_isFull;
    partialRound_tempInput_delay_46_payload_fullRound <= partialRound_tempInput_delay_45_payload_fullRound;
    partialRound_tempInput_delay_46_payload_partialRound <= partialRound_tempInput_delay_45_payload_partialRound;
    partialRound_tempInput_delay_46_payload_stateSize <= partialRound_tempInput_delay_45_payload_stateSize;
    partialRound_tempInput_delay_46_payload_stateID <= partialRound_tempInput_delay_45_payload_stateID;
    partialRound_tempInput_delay_46_payload_stateElements_0 <= partialRound_tempInput_delay_45_payload_stateElements_0;
    partialRound_tempInput_delay_46_payload_stateElements_1 <= partialRound_tempInput_delay_45_payload_stateElements_1;
    partialRound_tempInput_delay_46_payload_stateElements_2 <= partialRound_tempInput_delay_45_payload_stateElements_2;
    partialRound_tempInput_delay_46_payload_stateElements_3 <= partialRound_tempInput_delay_45_payload_stateElements_3;
    partialRound_tempInput_delay_46_payload_stateElements_4 <= partialRound_tempInput_delay_45_payload_stateElements_4;
    partialRound_tempInput_delay_46_payload_stateElements_5 <= partialRound_tempInput_delay_45_payload_stateElements_5;
    partialRound_tempInput_delay_46_payload_stateElements_6 <= partialRound_tempInput_delay_45_payload_stateElements_6;
    partialRound_tempInput_delay_46_payload_stateElements_7 <= partialRound_tempInput_delay_45_payload_stateElements_7;
    partialRound_tempInput_delay_46_payload_stateElements_8 <= partialRound_tempInput_delay_45_payload_stateElements_8;
    partialRound_tempInput_delay_46_payload_stateElements_9 <= partialRound_tempInput_delay_45_payload_stateElements_9;
    partialRound_tempInput_delay_46_payload_stateElements_10 <= partialRound_tempInput_delay_45_payload_stateElements_10;
    partialRound_tempInput_delay_46_payload_stateElements_11 <= partialRound_tempInput_delay_45_payload_stateElements_11;
    partialRound_tempInput_delay_47_valid <= partialRound_tempInput_delay_46_valid;
    partialRound_tempInput_delay_47_payload_isFull <= partialRound_tempInput_delay_46_payload_isFull;
    partialRound_tempInput_delay_47_payload_fullRound <= partialRound_tempInput_delay_46_payload_fullRound;
    partialRound_tempInput_delay_47_payload_partialRound <= partialRound_tempInput_delay_46_payload_partialRound;
    partialRound_tempInput_delay_47_payload_stateSize <= partialRound_tempInput_delay_46_payload_stateSize;
    partialRound_tempInput_delay_47_payload_stateID <= partialRound_tempInput_delay_46_payload_stateID;
    partialRound_tempInput_delay_47_payload_stateElements_0 <= partialRound_tempInput_delay_46_payload_stateElements_0;
    partialRound_tempInput_delay_47_payload_stateElements_1 <= partialRound_tempInput_delay_46_payload_stateElements_1;
    partialRound_tempInput_delay_47_payload_stateElements_2 <= partialRound_tempInput_delay_46_payload_stateElements_2;
    partialRound_tempInput_delay_47_payload_stateElements_3 <= partialRound_tempInput_delay_46_payload_stateElements_3;
    partialRound_tempInput_delay_47_payload_stateElements_4 <= partialRound_tempInput_delay_46_payload_stateElements_4;
    partialRound_tempInput_delay_47_payload_stateElements_5 <= partialRound_tempInput_delay_46_payload_stateElements_5;
    partialRound_tempInput_delay_47_payload_stateElements_6 <= partialRound_tempInput_delay_46_payload_stateElements_6;
    partialRound_tempInput_delay_47_payload_stateElements_7 <= partialRound_tempInput_delay_46_payload_stateElements_7;
    partialRound_tempInput_delay_47_payload_stateElements_8 <= partialRound_tempInput_delay_46_payload_stateElements_8;
    partialRound_tempInput_delay_47_payload_stateElements_9 <= partialRound_tempInput_delay_46_payload_stateElements_9;
    partialRound_tempInput_delay_47_payload_stateElements_10 <= partialRound_tempInput_delay_46_payload_stateElements_10;
    partialRound_tempInput_delay_47_payload_stateElements_11 <= partialRound_tempInput_delay_46_payload_stateElements_11;
    partialRound_tempInput_delay_48_valid <= partialRound_tempInput_delay_47_valid;
    partialRound_tempInput_delay_48_payload_isFull <= partialRound_tempInput_delay_47_payload_isFull;
    partialRound_tempInput_delay_48_payload_fullRound <= partialRound_tempInput_delay_47_payload_fullRound;
    partialRound_tempInput_delay_48_payload_partialRound <= partialRound_tempInput_delay_47_payload_partialRound;
    partialRound_tempInput_delay_48_payload_stateSize <= partialRound_tempInput_delay_47_payload_stateSize;
    partialRound_tempInput_delay_48_payload_stateID <= partialRound_tempInput_delay_47_payload_stateID;
    partialRound_tempInput_delay_48_payload_stateElements_0 <= partialRound_tempInput_delay_47_payload_stateElements_0;
    partialRound_tempInput_delay_48_payload_stateElements_1 <= partialRound_tempInput_delay_47_payload_stateElements_1;
    partialRound_tempInput_delay_48_payload_stateElements_2 <= partialRound_tempInput_delay_47_payload_stateElements_2;
    partialRound_tempInput_delay_48_payload_stateElements_3 <= partialRound_tempInput_delay_47_payload_stateElements_3;
    partialRound_tempInput_delay_48_payload_stateElements_4 <= partialRound_tempInput_delay_47_payload_stateElements_4;
    partialRound_tempInput_delay_48_payload_stateElements_5 <= partialRound_tempInput_delay_47_payload_stateElements_5;
    partialRound_tempInput_delay_48_payload_stateElements_6 <= partialRound_tempInput_delay_47_payload_stateElements_6;
    partialRound_tempInput_delay_48_payload_stateElements_7 <= partialRound_tempInput_delay_47_payload_stateElements_7;
    partialRound_tempInput_delay_48_payload_stateElements_8 <= partialRound_tempInput_delay_47_payload_stateElements_8;
    partialRound_tempInput_delay_48_payload_stateElements_9 <= partialRound_tempInput_delay_47_payload_stateElements_9;
    partialRound_tempInput_delay_48_payload_stateElements_10 <= partialRound_tempInput_delay_47_payload_stateElements_10;
    partialRound_tempInput_delay_48_payload_stateElements_11 <= partialRound_tempInput_delay_47_payload_stateElements_11;
    partialRound_tempInput_delay_49_valid <= partialRound_tempInput_delay_48_valid;
    partialRound_tempInput_delay_49_payload_isFull <= partialRound_tempInput_delay_48_payload_isFull;
    partialRound_tempInput_delay_49_payload_fullRound <= partialRound_tempInput_delay_48_payload_fullRound;
    partialRound_tempInput_delay_49_payload_partialRound <= partialRound_tempInput_delay_48_payload_partialRound;
    partialRound_tempInput_delay_49_payload_stateSize <= partialRound_tempInput_delay_48_payload_stateSize;
    partialRound_tempInput_delay_49_payload_stateID <= partialRound_tempInput_delay_48_payload_stateID;
    partialRound_tempInput_delay_49_payload_stateElements_0 <= partialRound_tempInput_delay_48_payload_stateElements_0;
    partialRound_tempInput_delay_49_payload_stateElements_1 <= partialRound_tempInput_delay_48_payload_stateElements_1;
    partialRound_tempInput_delay_49_payload_stateElements_2 <= partialRound_tempInput_delay_48_payload_stateElements_2;
    partialRound_tempInput_delay_49_payload_stateElements_3 <= partialRound_tempInput_delay_48_payload_stateElements_3;
    partialRound_tempInput_delay_49_payload_stateElements_4 <= partialRound_tempInput_delay_48_payload_stateElements_4;
    partialRound_tempInput_delay_49_payload_stateElements_5 <= partialRound_tempInput_delay_48_payload_stateElements_5;
    partialRound_tempInput_delay_49_payload_stateElements_6 <= partialRound_tempInput_delay_48_payload_stateElements_6;
    partialRound_tempInput_delay_49_payload_stateElements_7 <= partialRound_tempInput_delay_48_payload_stateElements_7;
    partialRound_tempInput_delay_49_payload_stateElements_8 <= partialRound_tempInput_delay_48_payload_stateElements_8;
    partialRound_tempInput_delay_49_payload_stateElements_9 <= partialRound_tempInput_delay_48_payload_stateElements_9;
    partialRound_tempInput_delay_49_payload_stateElements_10 <= partialRound_tempInput_delay_48_payload_stateElements_10;
    partialRound_tempInput_delay_49_payload_stateElements_11 <= partialRound_tempInput_delay_48_payload_stateElements_11;
    partialRound_tempInput_delay_50_valid <= partialRound_tempInput_delay_49_valid;
    partialRound_tempInput_delay_50_payload_isFull <= partialRound_tempInput_delay_49_payload_isFull;
    partialRound_tempInput_delay_50_payload_fullRound <= partialRound_tempInput_delay_49_payload_fullRound;
    partialRound_tempInput_delay_50_payload_partialRound <= partialRound_tempInput_delay_49_payload_partialRound;
    partialRound_tempInput_delay_50_payload_stateSize <= partialRound_tempInput_delay_49_payload_stateSize;
    partialRound_tempInput_delay_50_payload_stateID <= partialRound_tempInput_delay_49_payload_stateID;
    partialRound_tempInput_delay_50_payload_stateElements_0 <= partialRound_tempInput_delay_49_payload_stateElements_0;
    partialRound_tempInput_delay_50_payload_stateElements_1 <= partialRound_tempInput_delay_49_payload_stateElements_1;
    partialRound_tempInput_delay_50_payload_stateElements_2 <= partialRound_tempInput_delay_49_payload_stateElements_2;
    partialRound_tempInput_delay_50_payload_stateElements_3 <= partialRound_tempInput_delay_49_payload_stateElements_3;
    partialRound_tempInput_delay_50_payload_stateElements_4 <= partialRound_tempInput_delay_49_payload_stateElements_4;
    partialRound_tempInput_delay_50_payload_stateElements_5 <= partialRound_tempInput_delay_49_payload_stateElements_5;
    partialRound_tempInput_delay_50_payload_stateElements_6 <= partialRound_tempInput_delay_49_payload_stateElements_6;
    partialRound_tempInput_delay_50_payload_stateElements_7 <= partialRound_tempInput_delay_49_payload_stateElements_7;
    partialRound_tempInput_delay_50_payload_stateElements_8 <= partialRound_tempInput_delay_49_payload_stateElements_8;
    partialRound_tempInput_delay_50_payload_stateElements_9 <= partialRound_tempInput_delay_49_payload_stateElements_9;
    partialRound_tempInput_delay_50_payload_stateElements_10 <= partialRound_tempInput_delay_49_payload_stateElements_10;
    partialRound_tempInput_delay_50_payload_stateElements_11 <= partialRound_tempInput_delay_49_payload_stateElements_11;
    partialRound_tempInput_delay_51_valid <= partialRound_tempInput_delay_50_valid;
    partialRound_tempInput_delay_51_payload_isFull <= partialRound_tempInput_delay_50_payload_isFull;
    partialRound_tempInput_delay_51_payload_fullRound <= partialRound_tempInput_delay_50_payload_fullRound;
    partialRound_tempInput_delay_51_payload_partialRound <= partialRound_tempInput_delay_50_payload_partialRound;
    partialRound_tempInput_delay_51_payload_stateSize <= partialRound_tempInput_delay_50_payload_stateSize;
    partialRound_tempInput_delay_51_payload_stateID <= partialRound_tempInput_delay_50_payload_stateID;
    partialRound_tempInput_delay_51_payload_stateElements_0 <= partialRound_tempInput_delay_50_payload_stateElements_0;
    partialRound_tempInput_delay_51_payload_stateElements_1 <= partialRound_tempInput_delay_50_payload_stateElements_1;
    partialRound_tempInput_delay_51_payload_stateElements_2 <= partialRound_tempInput_delay_50_payload_stateElements_2;
    partialRound_tempInput_delay_51_payload_stateElements_3 <= partialRound_tempInput_delay_50_payload_stateElements_3;
    partialRound_tempInput_delay_51_payload_stateElements_4 <= partialRound_tempInput_delay_50_payload_stateElements_4;
    partialRound_tempInput_delay_51_payload_stateElements_5 <= partialRound_tempInput_delay_50_payload_stateElements_5;
    partialRound_tempInput_delay_51_payload_stateElements_6 <= partialRound_tempInput_delay_50_payload_stateElements_6;
    partialRound_tempInput_delay_51_payload_stateElements_7 <= partialRound_tempInput_delay_50_payload_stateElements_7;
    partialRound_tempInput_delay_51_payload_stateElements_8 <= partialRound_tempInput_delay_50_payload_stateElements_8;
    partialRound_tempInput_delay_51_payload_stateElements_9 <= partialRound_tempInput_delay_50_payload_stateElements_9;
    partialRound_tempInput_delay_51_payload_stateElements_10 <= partialRound_tempInput_delay_50_payload_stateElements_10;
    partialRound_tempInput_delay_51_payload_stateElements_11 <= partialRound_tempInput_delay_50_payload_stateElements_11;
    partialRound_tempInput_delay_52_valid <= partialRound_tempInput_delay_51_valid;
    partialRound_tempInput_delay_52_payload_isFull <= partialRound_tempInput_delay_51_payload_isFull;
    partialRound_tempInput_delay_52_payload_fullRound <= partialRound_tempInput_delay_51_payload_fullRound;
    partialRound_tempInput_delay_52_payload_partialRound <= partialRound_tempInput_delay_51_payload_partialRound;
    partialRound_tempInput_delay_52_payload_stateSize <= partialRound_tempInput_delay_51_payload_stateSize;
    partialRound_tempInput_delay_52_payload_stateID <= partialRound_tempInput_delay_51_payload_stateID;
    partialRound_tempInput_delay_52_payload_stateElements_0 <= partialRound_tempInput_delay_51_payload_stateElements_0;
    partialRound_tempInput_delay_52_payload_stateElements_1 <= partialRound_tempInput_delay_51_payload_stateElements_1;
    partialRound_tempInput_delay_52_payload_stateElements_2 <= partialRound_tempInput_delay_51_payload_stateElements_2;
    partialRound_tempInput_delay_52_payload_stateElements_3 <= partialRound_tempInput_delay_51_payload_stateElements_3;
    partialRound_tempInput_delay_52_payload_stateElements_4 <= partialRound_tempInput_delay_51_payload_stateElements_4;
    partialRound_tempInput_delay_52_payload_stateElements_5 <= partialRound_tempInput_delay_51_payload_stateElements_5;
    partialRound_tempInput_delay_52_payload_stateElements_6 <= partialRound_tempInput_delay_51_payload_stateElements_6;
    partialRound_tempInput_delay_52_payload_stateElements_7 <= partialRound_tempInput_delay_51_payload_stateElements_7;
    partialRound_tempInput_delay_52_payload_stateElements_8 <= partialRound_tempInput_delay_51_payload_stateElements_8;
    partialRound_tempInput_delay_52_payload_stateElements_9 <= partialRound_tempInput_delay_51_payload_stateElements_9;
    partialRound_tempInput_delay_52_payload_stateElements_10 <= partialRound_tempInput_delay_51_payload_stateElements_10;
    partialRound_tempInput_delay_52_payload_stateElements_11 <= partialRound_tempInput_delay_51_payload_stateElements_11;
    partialRound_tempInput_delay_53_valid <= partialRound_tempInput_delay_52_valid;
    partialRound_tempInput_delay_53_payload_isFull <= partialRound_tempInput_delay_52_payload_isFull;
    partialRound_tempInput_delay_53_payload_fullRound <= partialRound_tempInput_delay_52_payload_fullRound;
    partialRound_tempInput_delay_53_payload_partialRound <= partialRound_tempInput_delay_52_payload_partialRound;
    partialRound_tempInput_delay_53_payload_stateSize <= partialRound_tempInput_delay_52_payload_stateSize;
    partialRound_tempInput_delay_53_payload_stateID <= partialRound_tempInput_delay_52_payload_stateID;
    partialRound_tempInput_delay_53_payload_stateElements_0 <= partialRound_tempInput_delay_52_payload_stateElements_0;
    partialRound_tempInput_delay_53_payload_stateElements_1 <= partialRound_tempInput_delay_52_payload_stateElements_1;
    partialRound_tempInput_delay_53_payload_stateElements_2 <= partialRound_tempInput_delay_52_payload_stateElements_2;
    partialRound_tempInput_delay_53_payload_stateElements_3 <= partialRound_tempInput_delay_52_payload_stateElements_3;
    partialRound_tempInput_delay_53_payload_stateElements_4 <= partialRound_tempInput_delay_52_payload_stateElements_4;
    partialRound_tempInput_delay_53_payload_stateElements_5 <= partialRound_tempInput_delay_52_payload_stateElements_5;
    partialRound_tempInput_delay_53_payload_stateElements_6 <= partialRound_tempInput_delay_52_payload_stateElements_6;
    partialRound_tempInput_delay_53_payload_stateElements_7 <= partialRound_tempInput_delay_52_payload_stateElements_7;
    partialRound_tempInput_delay_53_payload_stateElements_8 <= partialRound_tempInput_delay_52_payload_stateElements_8;
    partialRound_tempInput_delay_53_payload_stateElements_9 <= partialRound_tempInput_delay_52_payload_stateElements_9;
    partialRound_tempInput_delay_53_payload_stateElements_10 <= partialRound_tempInput_delay_52_payload_stateElements_10;
    partialRound_tempInput_delay_53_payload_stateElements_11 <= partialRound_tempInput_delay_52_payload_stateElements_11;
    partialRound_tempInput_delay_54_valid <= partialRound_tempInput_delay_53_valid;
    partialRound_tempInput_delay_54_payload_isFull <= partialRound_tempInput_delay_53_payload_isFull;
    partialRound_tempInput_delay_54_payload_fullRound <= partialRound_tempInput_delay_53_payload_fullRound;
    partialRound_tempInput_delay_54_payload_partialRound <= partialRound_tempInput_delay_53_payload_partialRound;
    partialRound_tempInput_delay_54_payload_stateSize <= partialRound_tempInput_delay_53_payload_stateSize;
    partialRound_tempInput_delay_54_payload_stateID <= partialRound_tempInput_delay_53_payload_stateID;
    partialRound_tempInput_delay_54_payload_stateElements_0 <= partialRound_tempInput_delay_53_payload_stateElements_0;
    partialRound_tempInput_delay_54_payload_stateElements_1 <= partialRound_tempInput_delay_53_payload_stateElements_1;
    partialRound_tempInput_delay_54_payload_stateElements_2 <= partialRound_tempInput_delay_53_payload_stateElements_2;
    partialRound_tempInput_delay_54_payload_stateElements_3 <= partialRound_tempInput_delay_53_payload_stateElements_3;
    partialRound_tempInput_delay_54_payload_stateElements_4 <= partialRound_tempInput_delay_53_payload_stateElements_4;
    partialRound_tempInput_delay_54_payload_stateElements_5 <= partialRound_tempInput_delay_53_payload_stateElements_5;
    partialRound_tempInput_delay_54_payload_stateElements_6 <= partialRound_tempInput_delay_53_payload_stateElements_6;
    partialRound_tempInput_delay_54_payload_stateElements_7 <= partialRound_tempInput_delay_53_payload_stateElements_7;
    partialRound_tempInput_delay_54_payload_stateElements_8 <= partialRound_tempInput_delay_53_payload_stateElements_8;
    partialRound_tempInput_delay_54_payload_stateElements_9 <= partialRound_tempInput_delay_53_payload_stateElements_9;
    partialRound_tempInput_delay_54_payload_stateElements_10 <= partialRound_tempInput_delay_53_payload_stateElements_10;
    partialRound_tempInput_delay_54_payload_stateElements_11 <= partialRound_tempInput_delay_53_payload_stateElements_11;
    partialRound_tempInput_delay_55_valid <= partialRound_tempInput_delay_54_valid;
    partialRound_tempInput_delay_55_payload_isFull <= partialRound_tempInput_delay_54_payload_isFull;
    partialRound_tempInput_delay_55_payload_fullRound <= partialRound_tempInput_delay_54_payload_fullRound;
    partialRound_tempInput_delay_55_payload_partialRound <= partialRound_tempInput_delay_54_payload_partialRound;
    partialRound_tempInput_delay_55_payload_stateSize <= partialRound_tempInput_delay_54_payload_stateSize;
    partialRound_tempInput_delay_55_payload_stateID <= partialRound_tempInput_delay_54_payload_stateID;
    partialRound_tempInput_delay_55_payload_stateElements_0 <= partialRound_tempInput_delay_54_payload_stateElements_0;
    partialRound_tempInput_delay_55_payload_stateElements_1 <= partialRound_tempInput_delay_54_payload_stateElements_1;
    partialRound_tempInput_delay_55_payload_stateElements_2 <= partialRound_tempInput_delay_54_payload_stateElements_2;
    partialRound_tempInput_delay_55_payload_stateElements_3 <= partialRound_tempInput_delay_54_payload_stateElements_3;
    partialRound_tempInput_delay_55_payload_stateElements_4 <= partialRound_tempInput_delay_54_payload_stateElements_4;
    partialRound_tempInput_delay_55_payload_stateElements_5 <= partialRound_tempInput_delay_54_payload_stateElements_5;
    partialRound_tempInput_delay_55_payload_stateElements_6 <= partialRound_tempInput_delay_54_payload_stateElements_6;
    partialRound_tempInput_delay_55_payload_stateElements_7 <= partialRound_tempInput_delay_54_payload_stateElements_7;
    partialRound_tempInput_delay_55_payload_stateElements_8 <= partialRound_tempInput_delay_54_payload_stateElements_8;
    partialRound_tempInput_delay_55_payload_stateElements_9 <= partialRound_tempInput_delay_54_payload_stateElements_9;
    partialRound_tempInput_delay_55_payload_stateElements_10 <= partialRound_tempInput_delay_54_payload_stateElements_10;
    partialRound_tempInput_delay_55_payload_stateElements_11 <= partialRound_tempInput_delay_54_payload_stateElements_11;
    partialRound_tempInput_delay_56_valid <= partialRound_tempInput_delay_55_valid;
    partialRound_tempInput_delay_56_payload_isFull <= partialRound_tempInput_delay_55_payload_isFull;
    partialRound_tempInput_delay_56_payload_fullRound <= partialRound_tempInput_delay_55_payload_fullRound;
    partialRound_tempInput_delay_56_payload_partialRound <= partialRound_tempInput_delay_55_payload_partialRound;
    partialRound_tempInput_delay_56_payload_stateSize <= partialRound_tempInput_delay_55_payload_stateSize;
    partialRound_tempInput_delay_56_payload_stateID <= partialRound_tempInput_delay_55_payload_stateID;
    partialRound_tempInput_delay_56_payload_stateElements_0 <= partialRound_tempInput_delay_55_payload_stateElements_0;
    partialRound_tempInput_delay_56_payload_stateElements_1 <= partialRound_tempInput_delay_55_payload_stateElements_1;
    partialRound_tempInput_delay_56_payload_stateElements_2 <= partialRound_tempInput_delay_55_payload_stateElements_2;
    partialRound_tempInput_delay_56_payload_stateElements_3 <= partialRound_tempInput_delay_55_payload_stateElements_3;
    partialRound_tempInput_delay_56_payload_stateElements_4 <= partialRound_tempInput_delay_55_payload_stateElements_4;
    partialRound_tempInput_delay_56_payload_stateElements_5 <= partialRound_tempInput_delay_55_payload_stateElements_5;
    partialRound_tempInput_delay_56_payload_stateElements_6 <= partialRound_tempInput_delay_55_payload_stateElements_6;
    partialRound_tempInput_delay_56_payload_stateElements_7 <= partialRound_tempInput_delay_55_payload_stateElements_7;
    partialRound_tempInput_delay_56_payload_stateElements_8 <= partialRound_tempInput_delay_55_payload_stateElements_8;
    partialRound_tempInput_delay_56_payload_stateElements_9 <= partialRound_tempInput_delay_55_payload_stateElements_9;
    partialRound_tempInput_delay_56_payload_stateElements_10 <= partialRound_tempInput_delay_55_payload_stateElements_10;
    partialRound_tempInput_delay_56_payload_stateElements_11 <= partialRound_tempInput_delay_55_payload_stateElements_11;
    partialRound_tempInput_delay_57_valid <= partialRound_tempInput_delay_56_valid;
    partialRound_tempInput_delay_57_payload_isFull <= partialRound_tempInput_delay_56_payload_isFull;
    partialRound_tempInput_delay_57_payload_fullRound <= partialRound_tempInput_delay_56_payload_fullRound;
    partialRound_tempInput_delay_57_payload_partialRound <= partialRound_tempInput_delay_56_payload_partialRound;
    partialRound_tempInput_delay_57_payload_stateSize <= partialRound_tempInput_delay_56_payload_stateSize;
    partialRound_tempInput_delay_57_payload_stateID <= partialRound_tempInput_delay_56_payload_stateID;
    partialRound_tempInput_delay_57_payload_stateElements_0 <= partialRound_tempInput_delay_56_payload_stateElements_0;
    partialRound_tempInput_delay_57_payload_stateElements_1 <= partialRound_tempInput_delay_56_payload_stateElements_1;
    partialRound_tempInput_delay_57_payload_stateElements_2 <= partialRound_tempInput_delay_56_payload_stateElements_2;
    partialRound_tempInput_delay_57_payload_stateElements_3 <= partialRound_tempInput_delay_56_payload_stateElements_3;
    partialRound_tempInput_delay_57_payload_stateElements_4 <= partialRound_tempInput_delay_56_payload_stateElements_4;
    partialRound_tempInput_delay_57_payload_stateElements_5 <= partialRound_tempInput_delay_56_payload_stateElements_5;
    partialRound_tempInput_delay_57_payload_stateElements_6 <= partialRound_tempInput_delay_56_payload_stateElements_6;
    partialRound_tempInput_delay_57_payload_stateElements_7 <= partialRound_tempInput_delay_56_payload_stateElements_7;
    partialRound_tempInput_delay_57_payload_stateElements_8 <= partialRound_tempInput_delay_56_payload_stateElements_8;
    partialRound_tempInput_delay_57_payload_stateElements_9 <= partialRound_tempInput_delay_56_payload_stateElements_9;
    partialRound_tempInput_delay_57_payload_stateElements_10 <= partialRound_tempInput_delay_56_payload_stateElements_10;
    partialRound_tempInput_delay_57_payload_stateElements_11 <= partialRound_tempInput_delay_56_payload_stateElements_11;
    partialRound_tempInput_delay_58_valid <= partialRound_tempInput_delay_57_valid;
    partialRound_tempInput_delay_58_payload_isFull <= partialRound_tempInput_delay_57_payload_isFull;
    partialRound_tempInput_delay_58_payload_fullRound <= partialRound_tempInput_delay_57_payload_fullRound;
    partialRound_tempInput_delay_58_payload_partialRound <= partialRound_tempInput_delay_57_payload_partialRound;
    partialRound_tempInput_delay_58_payload_stateSize <= partialRound_tempInput_delay_57_payload_stateSize;
    partialRound_tempInput_delay_58_payload_stateID <= partialRound_tempInput_delay_57_payload_stateID;
    partialRound_tempInput_delay_58_payload_stateElements_0 <= partialRound_tempInput_delay_57_payload_stateElements_0;
    partialRound_tempInput_delay_58_payload_stateElements_1 <= partialRound_tempInput_delay_57_payload_stateElements_1;
    partialRound_tempInput_delay_58_payload_stateElements_2 <= partialRound_tempInput_delay_57_payload_stateElements_2;
    partialRound_tempInput_delay_58_payload_stateElements_3 <= partialRound_tempInput_delay_57_payload_stateElements_3;
    partialRound_tempInput_delay_58_payload_stateElements_4 <= partialRound_tempInput_delay_57_payload_stateElements_4;
    partialRound_tempInput_delay_58_payload_stateElements_5 <= partialRound_tempInput_delay_57_payload_stateElements_5;
    partialRound_tempInput_delay_58_payload_stateElements_6 <= partialRound_tempInput_delay_57_payload_stateElements_6;
    partialRound_tempInput_delay_58_payload_stateElements_7 <= partialRound_tempInput_delay_57_payload_stateElements_7;
    partialRound_tempInput_delay_58_payload_stateElements_8 <= partialRound_tempInput_delay_57_payload_stateElements_8;
    partialRound_tempInput_delay_58_payload_stateElements_9 <= partialRound_tempInput_delay_57_payload_stateElements_9;
    partialRound_tempInput_delay_58_payload_stateElements_10 <= partialRound_tempInput_delay_57_payload_stateElements_10;
    partialRound_tempInput_delay_58_payload_stateElements_11 <= partialRound_tempInput_delay_57_payload_stateElements_11;
    partialRound_tempInput_delay_59_valid <= partialRound_tempInput_delay_58_valid;
    partialRound_tempInput_delay_59_payload_isFull <= partialRound_tempInput_delay_58_payload_isFull;
    partialRound_tempInput_delay_59_payload_fullRound <= partialRound_tempInput_delay_58_payload_fullRound;
    partialRound_tempInput_delay_59_payload_partialRound <= partialRound_tempInput_delay_58_payload_partialRound;
    partialRound_tempInput_delay_59_payload_stateSize <= partialRound_tempInput_delay_58_payload_stateSize;
    partialRound_tempInput_delay_59_payload_stateID <= partialRound_tempInput_delay_58_payload_stateID;
    partialRound_tempInput_delay_59_payload_stateElements_0 <= partialRound_tempInput_delay_58_payload_stateElements_0;
    partialRound_tempInput_delay_59_payload_stateElements_1 <= partialRound_tempInput_delay_58_payload_stateElements_1;
    partialRound_tempInput_delay_59_payload_stateElements_2 <= partialRound_tempInput_delay_58_payload_stateElements_2;
    partialRound_tempInput_delay_59_payload_stateElements_3 <= partialRound_tempInput_delay_58_payload_stateElements_3;
    partialRound_tempInput_delay_59_payload_stateElements_4 <= partialRound_tempInput_delay_58_payload_stateElements_4;
    partialRound_tempInput_delay_59_payload_stateElements_5 <= partialRound_tempInput_delay_58_payload_stateElements_5;
    partialRound_tempInput_delay_59_payload_stateElements_6 <= partialRound_tempInput_delay_58_payload_stateElements_6;
    partialRound_tempInput_delay_59_payload_stateElements_7 <= partialRound_tempInput_delay_58_payload_stateElements_7;
    partialRound_tempInput_delay_59_payload_stateElements_8 <= partialRound_tempInput_delay_58_payload_stateElements_8;
    partialRound_tempInput_delay_59_payload_stateElements_9 <= partialRound_tempInput_delay_58_payload_stateElements_9;
    partialRound_tempInput_delay_59_payload_stateElements_10 <= partialRound_tempInput_delay_58_payload_stateElements_10;
    partialRound_tempInput_delay_59_payload_stateElements_11 <= partialRound_tempInput_delay_58_payload_stateElements_11;
    partialRound_tempInput_delay_60_valid <= partialRound_tempInput_delay_59_valid;
    partialRound_tempInput_delay_60_payload_isFull <= partialRound_tempInput_delay_59_payload_isFull;
    partialRound_tempInput_delay_60_payload_fullRound <= partialRound_tempInput_delay_59_payload_fullRound;
    partialRound_tempInput_delay_60_payload_partialRound <= partialRound_tempInput_delay_59_payload_partialRound;
    partialRound_tempInput_delay_60_payload_stateSize <= partialRound_tempInput_delay_59_payload_stateSize;
    partialRound_tempInput_delay_60_payload_stateID <= partialRound_tempInput_delay_59_payload_stateID;
    partialRound_tempInput_delay_60_payload_stateElements_0 <= partialRound_tempInput_delay_59_payload_stateElements_0;
    partialRound_tempInput_delay_60_payload_stateElements_1 <= partialRound_tempInput_delay_59_payload_stateElements_1;
    partialRound_tempInput_delay_60_payload_stateElements_2 <= partialRound_tempInput_delay_59_payload_stateElements_2;
    partialRound_tempInput_delay_60_payload_stateElements_3 <= partialRound_tempInput_delay_59_payload_stateElements_3;
    partialRound_tempInput_delay_60_payload_stateElements_4 <= partialRound_tempInput_delay_59_payload_stateElements_4;
    partialRound_tempInput_delay_60_payload_stateElements_5 <= partialRound_tempInput_delay_59_payload_stateElements_5;
    partialRound_tempInput_delay_60_payload_stateElements_6 <= partialRound_tempInput_delay_59_payload_stateElements_6;
    partialRound_tempInput_delay_60_payload_stateElements_7 <= partialRound_tempInput_delay_59_payload_stateElements_7;
    partialRound_tempInput_delay_60_payload_stateElements_8 <= partialRound_tempInput_delay_59_payload_stateElements_8;
    partialRound_tempInput_delay_60_payload_stateElements_9 <= partialRound_tempInput_delay_59_payload_stateElements_9;
    partialRound_tempInput_delay_60_payload_stateElements_10 <= partialRound_tempInput_delay_59_payload_stateElements_10;
    partialRound_tempInput_delay_60_payload_stateElements_11 <= partialRound_tempInput_delay_59_payload_stateElements_11;
    partialRound_tempInput_delay_61_valid <= partialRound_tempInput_delay_60_valid;
    partialRound_tempInput_delay_61_payload_isFull <= partialRound_tempInput_delay_60_payload_isFull;
    partialRound_tempInput_delay_61_payload_fullRound <= partialRound_tempInput_delay_60_payload_fullRound;
    partialRound_tempInput_delay_61_payload_partialRound <= partialRound_tempInput_delay_60_payload_partialRound;
    partialRound_tempInput_delay_61_payload_stateSize <= partialRound_tempInput_delay_60_payload_stateSize;
    partialRound_tempInput_delay_61_payload_stateID <= partialRound_tempInput_delay_60_payload_stateID;
    partialRound_tempInput_delay_61_payload_stateElements_0 <= partialRound_tempInput_delay_60_payload_stateElements_0;
    partialRound_tempInput_delay_61_payload_stateElements_1 <= partialRound_tempInput_delay_60_payload_stateElements_1;
    partialRound_tempInput_delay_61_payload_stateElements_2 <= partialRound_tempInput_delay_60_payload_stateElements_2;
    partialRound_tempInput_delay_61_payload_stateElements_3 <= partialRound_tempInput_delay_60_payload_stateElements_3;
    partialRound_tempInput_delay_61_payload_stateElements_4 <= partialRound_tempInput_delay_60_payload_stateElements_4;
    partialRound_tempInput_delay_61_payload_stateElements_5 <= partialRound_tempInput_delay_60_payload_stateElements_5;
    partialRound_tempInput_delay_61_payload_stateElements_6 <= partialRound_tempInput_delay_60_payload_stateElements_6;
    partialRound_tempInput_delay_61_payload_stateElements_7 <= partialRound_tempInput_delay_60_payload_stateElements_7;
    partialRound_tempInput_delay_61_payload_stateElements_8 <= partialRound_tempInput_delay_60_payload_stateElements_8;
    partialRound_tempInput_delay_61_payload_stateElements_9 <= partialRound_tempInput_delay_60_payload_stateElements_9;
    partialRound_tempInput_delay_61_payload_stateElements_10 <= partialRound_tempInput_delay_60_payload_stateElements_10;
    partialRound_tempInput_delay_61_payload_stateElements_11 <= partialRound_tempInput_delay_60_payload_stateElements_11;
    partialRound_tempInput_delay_62_valid <= partialRound_tempInput_delay_61_valid;
    partialRound_tempInput_delay_62_payload_isFull <= partialRound_tempInput_delay_61_payload_isFull;
    partialRound_tempInput_delay_62_payload_fullRound <= partialRound_tempInput_delay_61_payload_fullRound;
    partialRound_tempInput_delay_62_payload_partialRound <= partialRound_tempInput_delay_61_payload_partialRound;
    partialRound_tempInput_delay_62_payload_stateSize <= partialRound_tempInput_delay_61_payload_stateSize;
    partialRound_tempInput_delay_62_payload_stateID <= partialRound_tempInput_delay_61_payload_stateID;
    partialRound_tempInput_delay_62_payload_stateElements_0 <= partialRound_tempInput_delay_61_payload_stateElements_0;
    partialRound_tempInput_delay_62_payload_stateElements_1 <= partialRound_tempInput_delay_61_payload_stateElements_1;
    partialRound_tempInput_delay_62_payload_stateElements_2 <= partialRound_tempInput_delay_61_payload_stateElements_2;
    partialRound_tempInput_delay_62_payload_stateElements_3 <= partialRound_tempInput_delay_61_payload_stateElements_3;
    partialRound_tempInput_delay_62_payload_stateElements_4 <= partialRound_tempInput_delay_61_payload_stateElements_4;
    partialRound_tempInput_delay_62_payload_stateElements_5 <= partialRound_tempInput_delay_61_payload_stateElements_5;
    partialRound_tempInput_delay_62_payload_stateElements_6 <= partialRound_tempInput_delay_61_payload_stateElements_6;
    partialRound_tempInput_delay_62_payload_stateElements_7 <= partialRound_tempInput_delay_61_payload_stateElements_7;
    partialRound_tempInput_delay_62_payload_stateElements_8 <= partialRound_tempInput_delay_61_payload_stateElements_8;
    partialRound_tempInput_delay_62_payload_stateElements_9 <= partialRound_tempInput_delay_61_payload_stateElements_9;
    partialRound_tempInput_delay_62_payload_stateElements_10 <= partialRound_tempInput_delay_61_payload_stateElements_10;
    partialRound_tempInput_delay_62_payload_stateElements_11 <= partialRound_tempInput_delay_61_payload_stateElements_11;
    partialRound_tempInput_delay_63_valid <= partialRound_tempInput_delay_62_valid;
    partialRound_tempInput_delay_63_payload_isFull <= partialRound_tempInput_delay_62_payload_isFull;
    partialRound_tempInput_delay_63_payload_fullRound <= partialRound_tempInput_delay_62_payload_fullRound;
    partialRound_tempInput_delay_63_payload_partialRound <= partialRound_tempInput_delay_62_payload_partialRound;
    partialRound_tempInput_delay_63_payload_stateSize <= partialRound_tempInput_delay_62_payload_stateSize;
    partialRound_tempInput_delay_63_payload_stateID <= partialRound_tempInput_delay_62_payload_stateID;
    partialRound_tempInput_delay_63_payload_stateElements_0 <= partialRound_tempInput_delay_62_payload_stateElements_0;
    partialRound_tempInput_delay_63_payload_stateElements_1 <= partialRound_tempInput_delay_62_payload_stateElements_1;
    partialRound_tempInput_delay_63_payload_stateElements_2 <= partialRound_tempInput_delay_62_payload_stateElements_2;
    partialRound_tempInput_delay_63_payload_stateElements_3 <= partialRound_tempInput_delay_62_payload_stateElements_3;
    partialRound_tempInput_delay_63_payload_stateElements_4 <= partialRound_tempInput_delay_62_payload_stateElements_4;
    partialRound_tempInput_delay_63_payload_stateElements_5 <= partialRound_tempInput_delay_62_payload_stateElements_5;
    partialRound_tempInput_delay_63_payload_stateElements_6 <= partialRound_tempInput_delay_62_payload_stateElements_6;
    partialRound_tempInput_delay_63_payload_stateElements_7 <= partialRound_tempInput_delay_62_payload_stateElements_7;
    partialRound_tempInput_delay_63_payload_stateElements_8 <= partialRound_tempInput_delay_62_payload_stateElements_8;
    partialRound_tempInput_delay_63_payload_stateElements_9 <= partialRound_tempInput_delay_62_payload_stateElements_9;
    partialRound_tempInput_delay_63_payload_stateElements_10 <= partialRound_tempInput_delay_62_payload_stateElements_10;
    partialRound_tempInput_delay_63_payload_stateElements_11 <= partialRound_tempInput_delay_62_payload_stateElements_11;
    partialRound_contextDelayed_valid <= partialRound_tempInput_delay_63_valid;
    partialRound_contextDelayed_payload_isFull <= partialRound_tempInput_delay_63_payload_isFull;
    partialRound_contextDelayed_payload_fullRound <= partialRound_tempInput_delay_63_payload_fullRound;
    partialRound_contextDelayed_payload_partialRound <= partialRound_tempInput_delay_63_payload_partialRound;
    partialRound_contextDelayed_payload_stateSize <= partialRound_tempInput_delay_63_payload_stateSize;
    partialRound_contextDelayed_payload_stateID <= partialRound_tempInput_delay_63_payload_stateID;
    partialRound_contextDelayed_payload_stateElements_0 <= partialRound_tempInput_delay_63_payload_stateElements_0;
    partialRound_contextDelayed_payload_stateElements_1 <= partialRound_tempInput_delay_63_payload_stateElements_1;
    partialRound_contextDelayed_payload_stateElements_2 <= partialRound_tempInput_delay_63_payload_stateElements_2;
    partialRound_contextDelayed_payload_stateElements_3 <= partialRound_tempInput_delay_63_payload_stateElements_3;
    partialRound_contextDelayed_payload_stateElements_4 <= partialRound_tempInput_delay_63_payload_stateElements_4;
    partialRound_contextDelayed_payload_stateElements_5 <= partialRound_tempInput_delay_63_payload_stateElements_5;
    partialRound_contextDelayed_payload_stateElements_6 <= partialRound_tempInput_delay_63_payload_stateElements_6;
    partialRound_contextDelayed_payload_stateElements_7 <= partialRound_tempInput_delay_63_payload_stateElements_7;
    partialRound_contextDelayed_payload_stateElements_8 <= partialRound_tempInput_delay_63_payload_stateElements_8;
    partialRound_contextDelayed_payload_stateElements_9 <= partialRound_tempInput_delay_63_payload_stateElements_9;
    partialRound_contextDelayed_payload_stateElements_10 <= partialRound_tempInput_delay_63_payload_stateElements_10;
    partialRound_contextDelayed_payload_stateElements_11 <= partialRound_tempInput_delay_63_payload_stateElements_11;
    partialRound_output_payload_isFull <= partialRound_contextDelayed_payload_isFull;
    partialRound_output_payload_fullRound <= partialRound_contextDelayed_payload_fullRound;
    partialRound_output_payload_partialRound <= partialRound_contextDelayed_payload_partialRound;
    partialRound_output_payload_stateSize <= partialRound_contextDelayed_payload_stateSize;
    partialRound_output_payload_stateID <= partialRound_contextDelayed_payload_stateID;
    partialRound_output_payload_stateElements_0 <= _zz_partialRound_output_payload_stateElements_0;
    partialRound_output_payload_stateElements_1 <= partialRound_contextDelayed_payload_stateElements_1;
    partialRound_output_payload_stateElements_2 <= partialRound_contextDelayed_payload_stateElements_2;
    partialRound_output_payload_stateElements_3 <= _zz_partialRound_output_payload_stateElements_3;
    partialRound_output_payload_stateElements_4 <= _zz_partialRound_output_payload_stateElements_4;
    partialRound_output_payload_stateElements_5 <= _zz_partialRound_output_payload_stateElements_5;
    partialRound_output_payload_stateElements_6 <= _zz_partialRound_output_payload_stateElements_6;
    partialRound_output_payload_stateElements_7 <= _zz_partialRound_output_payload_stateElements_7;
    partialRound_output_payload_stateElements_8 <= _zz_partialRound_output_payload_stateElements_8;
    partialRound_output_payload_stateElements_9 <= partialRound_contextDelayed_payload_stateElements_9;
    partialRound_output_payload_stateElements_10 <= partialRound_contextDelayed_payload_stateElements_10;
    partialRound_output_payload_stateElements_11 <= partialRound_contextDelayed_payload_stateElements_11;
    fullRound_addContext_delay_1_valid <= fullRound_addContext_valid;
    fullRound_addContext_delay_1_payload_isFull <= fullRound_addContext_payload_isFull;
    fullRound_addContext_delay_1_payload_fullRound <= fullRound_addContext_payload_fullRound;
    fullRound_addContext_delay_1_payload_partialRound <= fullRound_addContext_payload_partialRound;
    fullRound_addContext_delay_1_payload_stateSize <= fullRound_addContext_payload_stateSize;
    fullRound_addContext_delay_1_payload_stateID <= fullRound_addContext_payload_stateID;
    fullRound_addContext_delay_2_valid <= fullRound_addContext_delay_1_valid;
    fullRound_addContext_delay_2_payload_isFull <= fullRound_addContext_delay_1_payload_isFull;
    fullRound_addContext_delay_2_payload_fullRound <= fullRound_addContext_delay_1_payload_fullRound;
    fullRound_addContext_delay_2_payload_partialRound <= fullRound_addContext_delay_1_payload_partialRound;
    fullRound_addContext_delay_2_payload_stateSize <= fullRound_addContext_delay_1_payload_stateSize;
    fullRound_addContext_delay_2_payload_stateID <= fullRound_addContext_delay_1_payload_stateID;
    fullRound_addContext_delay_3_valid <= fullRound_addContext_delay_2_valid;
    fullRound_addContext_delay_3_payload_isFull <= fullRound_addContext_delay_2_payload_isFull;
    fullRound_addContext_delay_3_payload_fullRound <= fullRound_addContext_delay_2_payload_fullRound;
    fullRound_addContext_delay_3_payload_partialRound <= fullRound_addContext_delay_2_payload_partialRound;
    fullRound_addContext_delay_3_payload_stateSize <= fullRound_addContext_delay_2_payload_stateSize;
    fullRound_addContext_delay_3_payload_stateID <= fullRound_addContext_delay_2_payload_stateID;
    fullRound_addContext_delay_4_valid <= fullRound_addContext_delay_3_valid;
    fullRound_addContext_delay_4_payload_isFull <= fullRound_addContext_delay_3_payload_isFull;
    fullRound_addContext_delay_4_payload_fullRound <= fullRound_addContext_delay_3_payload_fullRound;
    fullRound_addContext_delay_4_payload_partialRound <= fullRound_addContext_delay_3_payload_partialRound;
    fullRound_addContext_delay_4_payload_stateSize <= fullRound_addContext_delay_3_payload_stateSize;
    fullRound_addContext_delay_4_payload_stateID <= fullRound_addContext_delay_3_payload_stateID;
    fullRound_addContext_delay_5_valid <= fullRound_addContext_delay_4_valid;
    fullRound_addContext_delay_5_payload_isFull <= fullRound_addContext_delay_4_payload_isFull;
    fullRound_addContext_delay_5_payload_fullRound <= fullRound_addContext_delay_4_payload_fullRound;
    fullRound_addContext_delay_5_payload_partialRound <= fullRound_addContext_delay_4_payload_partialRound;
    fullRound_addContext_delay_5_payload_stateSize <= fullRound_addContext_delay_4_payload_stateSize;
    fullRound_addContext_delay_5_payload_stateID <= fullRound_addContext_delay_4_payload_stateID;
    fullRound_addContext_delay_6_valid <= fullRound_addContext_delay_5_valid;
    fullRound_addContext_delay_6_payload_isFull <= fullRound_addContext_delay_5_payload_isFull;
    fullRound_addContext_delay_6_payload_fullRound <= fullRound_addContext_delay_5_payload_fullRound;
    fullRound_addContext_delay_6_payload_partialRound <= fullRound_addContext_delay_5_payload_partialRound;
    fullRound_addContext_delay_6_payload_stateSize <= fullRound_addContext_delay_5_payload_stateSize;
    fullRound_addContext_delay_6_payload_stateID <= fullRound_addContext_delay_5_payload_stateID;
    fullRound_addContext_delay_7_valid <= fullRound_addContext_delay_6_valid;
    fullRound_addContext_delay_7_payload_isFull <= fullRound_addContext_delay_6_payload_isFull;
    fullRound_addContext_delay_7_payload_fullRound <= fullRound_addContext_delay_6_payload_fullRound;
    fullRound_addContext_delay_7_payload_partialRound <= fullRound_addContext_delay_6_payload_partialRound;
    fullRound_addContext_delay_7_payload_stateSize <= fullRound_addContext_delay_6_payload_stateSize;
    fullRound_addContext_delay_7_payload_stateID <= fullRound_addContext_delay_6_payload_stateID;
    fullRound_addContext_delay_8_valid <= fullRound_addContext_delay_7_valid;
    fullRound_addContext_delay_8_payload_isFull <= fullRound_addContext_delay_7_payload_isFull;
    fullRound_addContext_delay_8_payload_fullRound <= fullRound_addContext_delay_7_payload_fullRound;
    fullRound_addContext_delay_8_payload_partialRound <= fullRound_addContext_delay_7_payload_partialRound;
    fullRound_addContext_delay_8_payload_stateSize <= fullRound_addContext_delay_7_payload_stateSize;
    fullRound_addContext_delay_8_payload_stateID <= fullRound_addContext_delay_7_payload_stateID;
    fullRound_addContext_delay_9_valid <= fullRound_addContext_delay_8_valid;
    fullRound_addContext_delay_9_payload_isFull <= fullRound_addContext_delay_8_payload_isFull;
    fullRound_addContext_delay_9_payload_fullRound <= fullRound_addContext_delay_8_payload_fullRound;
    fullRound_addContext_delay_9_payload_partialRound <= fullRound_addContext_delay_8_payload_partialRound;
    fullRound_addContext_delay_9_payload_stateSize <= fullRound_addContext_delay_8_payload_stateSize;
    fullRound_addContext_delay_9_payload_stateID <= fullRound_addContext_delay_8_payload_stateID;
    fullRound_addContext_delay_10_valid <= fullRound_addContext_delay_9_valid;
    fullRound_addContext_delay_10_payload_isFull <= fullRound_addContext_delay_9_payload_isFull;
    fullRound_addContext_delay_10_payload_fullRound <= fullRound_addContext_delay_9_payload_fullRound;
    fullRound_addContext_delay_10_payload_partialRound <= fullRound_addContext_delay_9_payload_partialRound;
    fullRound_addContext_delay_10_payload_stateSize <= fullRound_addContext_delay_9_payload_stateSize;
    fullRound_addContext_delay_10_payload_stateID <= fullRound_addContext_delay_9_payload_stateID;
    fullRound_addContext_delay_11_valid <= fullRound_addContext_delay_10_valid;
    fullRound_addContext_delay_11_payload_isFull <= fullRound_addContext_delay_10_payload_isFull;
    fullRound_addContext_delay_11_payload_fullRound <= fullRound_addContext_delay_10_payload_fullRound;
    fullRound_addContext_delay_11_payload_partialRound <= fullRound_addContext_delay_10_payload_partialRound;
    fullRound_addContext_delay_11_payload_stateSize <= fullRound_addContext_delay_10_payload_stateSize;
    fullRound_addContext_delay_11_payload_stateID <= fullRound_addContext_delay_10_payload_stateID;
    fullRound_addContext_delay_12_valid <= fullRound_addContext_delay_11_valid;
    fullRound_addContext_delay_12_payload_isFull <= fullRound_addContext_delay_11_payload_isFull;
    fullRound_addContext_delay_12_payload_fullRound <= fullRound_addContext_delay_11_payload_fullRound;
    fullRound_addContext_delay_12_payload_partialRound <= fullRound_addContext_delay_11_payload_partialRound;
    fullRound_addContext_delay_12_payload_stateSize <= fullRound_addContext_delay_11_payload_stateSize;
    fullRound_addContext_delay_12_payload_stateID <= fullRound_addContext_delay_11_payload_stateID;
    fullRound_addContext_delay_13_valid <= fullRound_addContext_delay_12_valid;
    fullRound_addContext_delay_13_payload_isFull <= fullRound_addContext_delay_12_payload_isFull;
    fullRound_addContext_delay_13_payload_fullRound <= fullRound_addContext_delay_12_payload_fullRound;
    fullRound_addContext_delay_13_payload_partialRound <= fullRound_addContext_delay_12_payload_partialRound;
    fullRound_addContext_delay_13_payload_stateSize <= fullRound_addContext_delay_12_payload_stateSize;
    fullRound_addContext_delay_13_payload_stateID <= fullRound_addContext_delay_12_payload_stateID;
    fullRound_addContext_delay_14_valid <= fullRound_addContext_delay_13_valid;
    fullRound_addContext_delay_14_payload_isFull <= fullRound_addContext_delay_13_payload_isFull;
    fullRound_addContext_delay_14_payload_fullRound <= fullRound_addContext_delay_13_payload_fullRound;
    fullRound_addContext_delay_14_payload_partialRound <= fullRound_addContext_delay_13_payload_partialRound;
    fullRound_addContext_delay_14_payload_stateSize <= fullRound_addContext_delay_13_payload_stateSize;
    fullRound_addContext_delay_14_payload_stateID <= fullRound_addContext_delay_13_payload_stateID;
    fullRound_addContext_delay_15_valid <= fullRound_addContext_delay_14_valid;
    fullRound_addContext_delay_15_payload_isFull <= fullRound_addContext_delay_14_payload_isFull;
    fullRound_addContext_delay_15_payload_fullRound <= fullRound_addContext_delay_14_payload_fullRound;
    fullRound_addContext_delay_15_payload_partialRound <= fullRound_addContext_delay_14_payload_partialRound;
    fullRound_addContext_delay_15_payload_stateSize <= fullRound_addContext_delay_14_payload_stateSize;
    fullRound_addContext_delay_15_payload_stateID <= fullRound_addContext_delay_14_payload_stateID;
    fullRound_addContext_delay_16_valid <= fullRound_addContext_delay_15_valid;
    fullRound_addContext_delay_16_payload_isFull <= fullRound_addContext_delay_15_payload_isFull;
    fullRound_addContext_delay_16_payload_fullRound <= fullRound_addContext_delay_15_payload_fullRound;
    fullRound_addContext_delay_16_payload_partialRound <= fullRound_addContext_delay_15_payload_partialRound;
    fullRound_addContext_delay_16_payload_stateSize <= fullRound_addContext_delay_15_payload_stateSize;
    fullRound_addContext_delay_16_payload_stateID <= fullRound_addContext_delay_15_payload_stateID;
    fullRound_addContext_delay_17_valid <= fullRound_addContext_delay_16_valid;
    fullRound_addContext_delay_17_payload_isFull <= fullRound_addContext_delay_16_payload_isFull;
    fullRound_addContext_delay_17_payload_fullRound <= fullRound_addContext_delay_16_payload_fullRound;
    fullRound_addContext_delay_17_payload_partialRound <= fullRound_addContext_delay_16_payload_partialRound;
    fullRound_addContext_delay_17_payload_stateSize <= fullRound_addContext_delay_16_payload_stateSize;
    fullRound_addContext_delay_17_payload_stateID <= fullRound_addContext_delay_16_payload_stateID;
    fullRound_addContext_delay_18_valid <= fullRound_addContext_delay_17_valid;
    fullRound_addContext_delay_18_payload_isFull <= fullRound_addContext_delay_17_payload_isFull;
    fullRound_addContext_delay_18_payload_fullRound <= fullRound_addContext_delay_17_payload_fullRound;
    fullRound_addContext_delay_18_payload_partialRound <= fullRound_addContext_delay_17_payload_partialRound;
    fullRound_addContext_delay_18_payload_stateSize <= fullRound_addContext_delay_17_payload_stateSize;
    fullRound_addContext_delay_18_payload_stateID <= fullRound_addContext_delay_17_payload_stateID;
    fullRound_addContext_delay_19_valid <= fullRound_addContext_delay_18_valid;
    fullRound_addContext_delay_19_payload_isFull <= fullRound_addContext_delay_18_payload_isFull;
    fullRound_addContext_delay_19_payload_fullRound <= fullRound_addContext_delay_18_payload_fullRound;
    fullRound_addContext_delay_19_payload_partialRound <= fullRound_addContext_delay_18_payload_partialRound;
    fullRound_addContext_delay_19_payload_stateSize <= fullRound_addContext_delay_18_payload_stateSize;
    fullRound_addContext_delay_19_payload_stateID <= fullRound_addContext_delay_18_payload_stateID;
    fullRound_addContext_delay_20_valid <= fullRound_addContext_delay_19_valid;
    fullRound_addContext_delay_20_payload_isFull <= fullRound_addContext_delay_19_payload_isFull;
    fullRound_addContext_delay_20_payload_fullRound <= fullRound_addContext_delay_19_payload_fullRound;
    fullRound_addContext_delay_20_payload_partialRound <= fullRound_addContext_delay_19_payload_partialRound;
    fullRound_addContext_delay_20_payload_stateSize <= fullRound_addContext_delay_19_payload_stateSize;
    fullRound_addContext_delay_20_payload_stateID <= fullRound_addContext_delay_19_payload_stateID;
    fullRound_addContext_delay_21_valid <= fullRound_addContext_delay_20_valid;
    fullRound_addContext_delay_21_payload_isFull <= fullRound_addContext_delay_20_payload_isFull;
    fullRound_addContext_delay_21_payload_fullRound <= fullRound_addContext_delay_20_payload_fullRound;
    fullRound_addContext_delay_21_payload_partialRound <= fullRound_addContext_delay_20_payload_partialRound;
    fullRound_addContext_delay_21_payload_stateSize <= fullRound_addContext_delay_20_payload_stateSize;
    fullRound_addContext_delay_21_payload_stateID <= fullRound_addContext_delay_20_payload_stateID;
    fullRound_addContext_delay_22_valid <= fullRound_addContext_delay_21_valid;
    fullRound_addContext_delay_22_payload_isFull <= fullRound_addContext_delay_21_payload_isFull;
    fullRound_addContext_delay_22_payload_fullRound <= fullRound_addContext_delay_21_payload_fullRound;
    fullRound_addContext_delay_22_payload_partialRound <= fullRound_addContext_delay_21_payload_partialRound;
    fullRound_addContext_delay_22_payload_stateSize <= fullRound_addContext_delay_21_payload_stateSize;
    fullRound_addContext_delay_22_payload_stateID <= fullRound_addContext_delay_21_payload_stateID;
    fullRound_addContext_delay_23_valid <= fullRound_addContext_delay_22_valid;
    fullRound_addContext_delay_23_payload_isFull <= fullRound_addContext_delay_22_payload_isFull;
    fullRound_addContext_delay_23_payload_fullRound <= fullRound_addContext_delay_22_payload_fullRound;
    fullRound_addContext_delay_23_payload_partialRound <= fullRound_addContext_delay_22_payload_partialRound;
    fullRound_addContext_delay_23_payload_stateSize <= fullRound_addContext_delay_22_payload_stateSize;
    fullRound_addContext_delay_23_payload_stateID <= fullRound_addContext_delay_22_payload_stateID;
    fullRound_addContext_delay_24_valid <= fullRound_addContext_delay_23_valid;
    fullRound_addContext_delay_24_payload_isFull <= fullRound_addContext_delay_23_payload_isFull;
    fullRound_addContext_delay_24_payload_fullRound <= fullRound_addContext_delay_23_payload_fullRound;
    fullRound_addContext_delay_24_payload_partialRound <= fullRound_addContext_delay_23_payload_partialRound;
    fullRound_addContext_delay_24_payload_stateSize <= fullRound_addContext_delay_23_payload_stateSize;
    fullRound_addContext_delay_24_payload_stateID <= fullRound_addContext_delay_23_payload_stateID;
    fullRound_addContext_delay_25_valid <= fullRound_addContext_delay_24_valid;
    fullRound_addContext_delay_25_payload_isFull <= fullRound_addContext_delay_24_payload_isFull;
    fullRound_addContext_delay_25_payload_fullRound <= fullRound_addContext_delay_24_payload_fullRound;
    fullRound_addContext_delay_25_payload_partialRound <= fullRound_addContext_delay_24_payload_partialRound;
    fullRound_addContext_delay_25_payload_stateSize <= fullRound_addContext_delay_24_payload_stateSize;
    fullRound_addContext_delay_25_payload_stateID <= fullRound_addContext_delay_24_payload_stateID;
    fullRound_addContext_delay_26_valid <= fullRound_addContext_delay_25_valid;
    fullRound_addContext_delay_26_payload_isFull <= fullRound_addContext_delay_25_payload_isFull;
    fullRound_addContext_delay_26_payload_fullRound <= fullRound_addContext_delay_25_payload_fullRound;
    fullRound_addContext_delay_26_payload_partialRound <= fullRound_addContext_delay_25_payload_partialRound;
    fullRound_addContext_delay_26_payload_stateSize <= fullRound_addContext_delay_25_payload_stateSize;
    fullRound_addContext_delay_26_payload_stateID <= fullRound_addContext_delay_25_payload_stateID;
    fullRound_addContext_delay_27_valid <= fullRound_addContext_delay_26_valid;
    fullRound_addContext_delay_27_payload_isFull <= fullRound_addContext_delay_26_payload_isFull;
    fullRound_addContext_delay_27_payload_fullRound <= fullRound_addContext_delay_26_payload_fullRound;
    fullRound_addContext_delay_27_payload_partialRound <= fullRound_addContext_delay_26_payload_partialRound;
    fullRound_addContext_delay_27_payload_stateSize <= fullRound_addContext_delay_26_payload_stateSize;
    fullRound_addContext_delay_27_payload_stateID <= fullRound_addContext_delay_26_payload_stateID;
    fullRound_addContext_delay_28_valid <= fullRound_addContext_delay_27_valid;
    fullRound_addContext_delay_28_payload_isFull <= fullRound_addContext_delay_27_payload_isFull;
    fullRound_addContext_delay_28_payload_fullRound <= fullRound_addContext_delay_27_payload_fullRound;
    fullRound_addContext_delay_28_payload_partialRound <= fullRound_addContext_delay_27_payload_partialRound;
    fullRound_addContext_delay_28_payload_stateSize <= fullRound_addContext_delay_27_payload_stateSize;
    fullRound_addContext_delay_28_payload_stateID <= fullRound_addContext_delay_27_payload_stateID;
    fullRound_addContext_delay_29_valid <= fullRound_addContext_delay_28_valid;
    fullRound_addContext_delay_29_payload_isFull <= fullRound_addContext_delay_28_payload_isFull;
    fullRound_addContext_delay_29_payload_fullRound <= fullRound_addContext_delay_28_payload_fullRound;
    fullRound_addContext_delay_29_payload_partialRound <= fullRound_addContext_delay_28_payload_partialRound;
    fullRound_addContext_delay_29_payload_stateSize <= fullRound_addContext_delay_28_payload_stateSize;
    fullRound_addContext_delay_29_payload_stateID <= fullRound_addContext_delay_28_payload_stateID;
    fullRound_addContext_delay_30_valid <= fullRound_addContext_delay_29_valid;
    fullRound_addContext_delay_30_payload_isFull <= fullRound_addContext_delay_29_payload_isFull;
    fullRound_addContext_delay_30_payload_fullRound <= fullRound_addContext_delay_29_payload_fullRound;
    fullRound_addContext_delay_30_payload_partialRound <= fullRound_addContext_delay_29_payload_partialRound;
    fullRound_addContext_delay_30_payload_stateSize <= fullRound_addContext_delay_29_payload_stateSize;
    fullRound_addContext_delay_30_payload_stateID <= fullRound_addContext_delay_29_payload_stateID;
    fullRound_addContext_delay_31_valid <= fullRound_addContext_delay_30_valid;
    fullRound_addContext_delay_31_payload_isFull <= fullRound_addContext_delay_30_payload_isFull;
    fullRound_addContext_delay_31_payload_fullRound <= fullRound_addContext_delay_30_payload_fullRound;
    fullRound_addContext_delay_31_payload_partialRound <= fullRound_addContext_delay_30_payload_partialRound;
    fullRound_addContext_delay_31_payload_stateSize <= fullRound_addContext_delay_30_payload_stateSize;
    fullRound_addContext_delay_31_payload_stateID <= fullRound_addContext_delay_30_payload_stateID;
    fullRound_addContext_delay_32_valid <= fullRound_addContext_delay_31_valid;
    fullRound_addContext_delay_32_payload_isFull <= fullRound_addContext_delay_31_payload_isFull;
    fullRound_addContext_delay_32_payload_fullRound <= fullRound_addContext_delay_31_payload_fullRound;
    fullRound_addContext_delay_32_payload_partialRound <= fullRound_addContext_delay_31_payload_partialRound;
    fullRound_addContext_delay_32_payload_stateSize <= fullRound_addContext_delay_31_payload_stateSize;
    fullRound_addContext_delay_32_payload_stateID <= fullRound_addContext_delay_31_payload_stateID;
    fullRound_addContext_delay_33_valid <= fullRound_addContext_delay_32_valid;
    fullRound_addContext_delay_33_payload_isFull <= fullRound_addContext_delay_32_payload_isFull;
    fullRound_addContext_delay_33_payload_fullRound <= fullRound_addContext_delay_32_payload_fullRound;
    fullRound_addContext_delay_33_payload_partialRound <= fullRound_addContext_delay_32_payload_partialRound;
    fullRound_addContext_delay_33_payload_stateSize <= fullRound_addContext_delay_32_payload_stateSize;
    fullRound_addContext_delay_33_payload_stateID <= fullRound_addContext_delay_32_payload_stateID;
    fullRound_addContext_delay_34_valid <= fullRound_addContext_delay_33_valid;
    fullRound_addContext_delay_34_payload_isFull <= fullRound_addContext_delay_33_payload_isFull;
    fullRound_addContext_delay_34_payload_fullRound <= fullRound_addContext_delay_33_payload_fullRound;
    fullRound_addContext_delay_34_payload_partialRound <= fullRound_addContext_delay_33_payload_partialRound;
    fullRound_addContext_delay_34_payload_stateSize <= fullRound_addContext_delay_33_payload_stateSize;
    fullRound_addContext_delay_34_payload_stateID <= fullRound_addContext_delay_33_payload_stateID;
    fullRound_addContext_delay_35_valid <= fullRound_addContext_delay_34_valid;
    fullRound_addContext_delay_35_payload_isFull <= fullRound_addContext_delay_34_payload_isFull;
    fullRound_addContext_delay_35_payload_fullRound <= fullRound_addContext_delay_34_payload_fullRound;
    fullRound_addContext_delay_35_payload_partialRound <= fullRound_addContext_delay_34_payload_partialRound;
    fullRound_addContext_delay_35_payload_stateSize <= fullRound_addContext_delay_34_payload_stateSize;
    fullRound_addContext_delay_35_payload_stateID <= fullRound_addContext_delay_34_payload_stateID;
    fullRound_addContext_delay_36_valid <= fullRound_addContext_delay_35_valid;
    fullRound_addContext_delay_36_payload_isFull <= fullRound_addContext_delay_35_payload_isFull;
    fullRound_addContext_delay_36_payload_fullRound <= fullRound_addContext_delay_35_payload_fullRound;
    fullRound_addContext_delay_36_payload_partialRound <= fullRound_addContext_delay_35_payload_partialRound;
    fullRound_addContext_delay_36_payload_stateSize <= fullRound_addContext_delay_35_payload_stateSize;
    fullRound_addContext_delay_36_payload_stateID <= fullRound_addContext_delay_35_payload_stateID;
    fullRound_addContext_delay_37_valid <= fullRound_addContext_delay_36_valid;
    fullRound_addContext_delay_37_payload_isFull <= fullRound_addContext_delay_36_payload_isFull;
    fullRound_addContext_delay_37_payload_fullRound <= fullRound_addContext_delay_36_payload_fullRound;
    fullRound_addContext_delay_37_payload_partialRound <= fullRound_addContext_delay_36_payload_partialRound;
    fullRound_addContext_delay_37_payload_stateSize <= fullRound_addContext_delay_36_payload_stateSize;
    fullRound_addContext_delay_37_payload_stateID <= fullRound_addContext_delay_36_payload_stateID;
    fullRound_addContext_delay_38_valid <= fullRound_addContext_delay_37_valid;
    fullRound_addContext_delay_38_payload_isFull <= fullRound_addContext_delay_37_payload_isFull;
    fullRound_addContext_delay_38_payload_fullRound <= fullRound_addContext_delay_37_payload_fullRound;
    fullRound_addContext_delay_38_payload_partialRound <= fullRound_addContext_delay_37_payload_partialRound;
    fullRound_addContext_delay_38_payload_stateSize <= fullRound_addContext_delay_37_payload_stateSize;
    fullRound_addContext_delay_38_payload_stateID <= fullRound_addContext_delay_37_payload_stateID;
    fullRound_addContext_delay_39_valid <= fullRound_addContext_delay_38_valid;
    fullRound_addContext_delay_39_payload_isFull <= fullRound_addContext_delay_38_payload_isFull;
    fullRound_addContext_delay_39_payload_fullRound <= fullRound_addContext_delay_38_payload_fullRound;
    fullRound_addContext_delay_39_payload_partialRound <= fullRound_addContext_delay_38_payload_partialRound;
    fullRound_addContext_delay_39_payload_stateSize <= fullRound_addContext_delay_38_payload_stateSize;
    fullRound_addContext_delay_39_payload_stateID <= fullRound_addContext_delay_38_payload_stateID;
    fullRound_addContext_delay_40_valid <= fullRound_addContext_delay_39_valid;
    fullRound_addContext_delay_40_payload_isFull <= fullRound_addContext_delay_39_payload_isFull;
    fullRound_addContext_delay_40_payload_fullRound <= fullRound_addContext_delay_39_payload_fullRound;
    fullRound_addContext_delay_40_payload_partialRound <= fullRound_addContext_delay_39_payload_partialRound;
    fullRound_addContext_delay_40_payload_stateSize <= fullRound_addContext_delay_39_payload_stateSize;
    fullRound_addContext_delay_40_payload_stateID <= fullRound_addContext_delay_39_payload_stateID;
    fullRound_addContext_delay_41_valid <= fullRound_addContext_delay_40_valid;
    fullRound_addContext_delay_41_payload_isFull <= fullRound_addContext_delay_40_payload_isFull;
    fullRound_addContext_delay_41_payload_fullRound <= fullRound_addContext_delay_40_payload_fullRound;
    fullRound_addContext_delay_41_payload_partialRound <= fullRound_addContext_delay_40_payload_partialRound;
    fullRound_addContext_delay_41_payload_stateSize <= fullRound_addContext_delay_40_payload_stateSize;
    fullRound_addContext_delay_41_payload_stateID <= fullRound_addContext_delay_40_payload_stateID;
    fullRound_addContext_delay_42_valid <= fullRound_addContext_delay_41_valid;
    fullRound_addContext_delay_42_payload_isFull <= fullRound_addContext_delay_41_payload_isFull;
    fullRound_addContext_delay_42_payload_fullRound <= fullRound_addContext_delay_41_payload_fullRound;
    fullRound_addContext_delay_42_payload_partialRound <= fullRound_addContext_delay_41_payload_partialRound;
    fullRound_addContext_delay_42_payload_stateSize <= fullRound_addContext_delay_41_payload_stateSize;
    fullRound_addContext_delay_42_payload_stateID <= fullRound_addContext_delay_41_payload_stateID;
    fullRound_addContext_delay_43_valid <= fullRound_addContext_delay_42_valid;
    fullRound_addContext_delay_43_payload_isFull <= fullRound_addContext_delay_42_payload_isFull;
    fullRound_addContext_delay_43_payload_fullRound <= fullRound_addContext_delay_42_payload_fullRound;
    fullRound_addContext_delay_43_payload_partialRound <= fullRound_addContext_delay_42_payload_partialRound;
    fullRound_addContext_delay_43_payload_stateSize <= fullRound_addContext_delay_42_payload_stateSize;
    fullRound_addContext_delay_43_payload_stateID <= fullRound_addContext_delay_42_payload_stateID;
    fullRound_addContext_delay_44_valid <= fullRound_addContext_delay_43_valid;
    fullRound_addContext_delay_44_payload_isFull <= fullRound_addContext_delay_43_payload_isFull;
    fullRound_addContext_delay_44_payload_fullRound <= fullRound_addContext_delay_43_payload_fullRound;
    fullRound_addContext_delay_44_payload_partialRound <= fullRound_addContext_delay_43_payload_partialRound;
    fullRound_addContext_delay_44_payload_stateSize <= fullRound_addContext_delay_43_payload_stateSize;
    fullRound_addContext_delay_44_payload_stateID <= fullRound_addContext_delay_43_payload_stateID;
    fullRound_addContext_delay_45_valid <= fullRound_addContext_delay_44_valid;
    fullRound_addContext_delay_45_payload_isFull <= fullRound_addContext_delay_44_payload_isFull;
    fullRound_addContext_delay_45_payload_fullRound <= fullRound_addContext_delay_44_payload_fullRound;
    fullRound_addContext_delay_45_payload_partialRound <= fullRound_addContext_delay_44_payload_partialRound;
    fullRound_addContext_delay_45_payload_stateSize <= fullRound_addContext_delay_44_payload_stateSize;
    fullRound_addContext_delay_45_payload_stateID <= fullRound_addContext_delay_44_payload_stateID;
    fullRound_addContext_delay_46_valid <= fullRound_addContext_delay_45_valid;
    fullRound_addContext_delay_46_payload_isFull <= fullRound_addContext_delay_45_payload_isFull;
    fullRound_addContext_delay_46_payload_fullRound <= fullRound_addContext_delay_45_payload_fullRound;
    fullRound_addContext_delay_46_payload_partialRound <= fullRound_addContext_delay_45_payload_partialRound;
    fullRound_addContext_delay_46_payload_stateSize <= fullRound_addContext_delay_45_payload_stateSize;
    fullRound_addContext_delay_46_payload_stateID <= fullRound_addContext_delay_45_payload_stateID;
    fullRound_addContext_delay_47_valid <= fullRound_addContext_delay_46_valid;
    fullRound_addContext_delay_47_payload_isFull <= fullRound_addContext_delay_46_payload_isFull;
    fullRound_addContext_delay_47_payload_fullRound <= fullRound_addContext_delay_46_payload_fullRound;
    fullRound_addContext_delay_47_payload_partialRound <= fullRound_addContext_delay_46_payload_partialRound;
    fullRound_addContext_delay_47_payload_stateSize <= fullRound_addContext_delay_46_payload_stateSize;
    fullRound_addContext_delay_47_payload_stateID <= fullRound_addContext_delay_46_payload_stateID;
    fullRound_addContext_delay_48_valid <= fullRound_addContext_delay_47_valid;
    fullRound_addContext_delay_48_payload_isFull <= fullRound_addContext_delay_47_payload_isFull;
    fullRound_addContext_delay_48_payload_fullRound <= fullRound_addContext_delay_47_payload_fullRound;
    fullRound_addContext_delay_48_payload_partialRound <= fullRound_addContext_delay_47_payload_partialRound;
    fullRound_addContext_delay_48_payload_stateSize <= fullRound_addContext_delay_47_payload_stateSize;
    fullRound_addContext_delay_48_payload_stateID <= fullRound_addContext_delay_47_payload_stateID;
    fullRound_addContext_delay_49_valid <= fullRound_addContext_delay_48_valid;
    fullRound_addContext_delay_49_payload_isFull <= fullRound_addContext_delay_48_payload_isFull;
    fullRound_addContext_delay_49_payload_fullRound <= fullRound_addContext_delay_48_payload_fullRound;
    fullRound_addContext_delay_49_payload_partialRound <= fullRound_addContext_delay_48_payload_partialRound;
    fullRound_addContext_delay_49_payload_stateSize <= fullRound_addContext_delay_48_payload_stateSize;
    fullRound_addContext_delay_49_payload_stateID <= fullRound_addContext_delay_48_payload_stateID;
    fullRound_addContext_delay_50_valid <= fullRound_addContext_delay_49_valid;
    fullRound_addContext_delay_50_payload_isFull <= fullRound_addContext_delay_49_payload_isFull;
    fullRound_addContext_delay_50_payload_fullRound <= fullRound_addContext_delay_49_payload_fullRound;
    fullRound_addContext_delay_50_payload_partialRound <= fullRound_addContext_delay_49_payload_partialRound;
    fullRound_addContext_delay_50_payload_stateSize <= fullRound_addContext_delay_49_payload_stateSize;
    fullRound_addContext_delay_50_payload_stateID <= fullRound_addContext_delay_49_payload_stateID;
    fullRound_addContext_delay_51_valid <= fullRound_addContext_delay_50_valid;
    fullRound_addContext_delay_51_payload_isFull <= fullRound_addContext_delay_50_payload_isFull;
    fullRound_addContext_delay_51_payload_fullRound <= fullRound_addContext_delay_50_payload_fullRound;
    fullRound_addContext_delay_51_payload_partialRound <= fullRound_addContext_delay_50_payload_partialRound;
    fullRound_addContext_delay_51_payload_stateSize <= fullRound_addContext_delay_50_payload_stateSize;
    fullRound_addContext_delay_51_payload_stateID <= fullRound_addContext_delay_50_payload_stateID;
    fullRound_addContext_delay_52_valid <= fullRound_addContext_delay_51_valid;
    fullRound_addContext_delay_52_payload_isFull <= fullRound_addContext_delay_51_payload_isFull;
    fullRound_addContext_delay_52_payload_fullRound <= fullRound_addContext_delay_51_payload_fullRound;
    fullRound_addContext_delay_52_payload_partialRound <= fullRound_addContext_delay_51_payload_partialRound;
    fullRound_addContext_delay_52_payload_stateSize <= fullRound_addContext_delay_51_payload_stateSize;
    fullRound_addContext_delay_52_payload_stateID <= fullRound_addContext_delay_51_payload_stateID;
    fullRound_addContext_delay_53_valid <= fullRound_addContext_delay_52_valid;
    fullRound_addContext_delay_53_payload_isFull <= fullRound_addContext_delay_52_payload_isFull;
    fullRound_addContext_delay_53_payload_fullRound <= fullRound_addContext_delay_52_payload_fullRound;
    fullRound_addContext_delay_53_payload_partialRound <= fullRound_addContext_delay_52_payload_partialRound;
    fullRound_addContext_delay_53_payload_stateSize <= fullRound_addContext_delay_52_payload_stateSize;
    fullRound_addContext_delay_53_payload_stateID <= fullRound_addContext_delay_52_payload_stateID;
    fullRound_addContext_delay_54_valid <= fullRound_addContext_delay_53_valid;
    fullRound_addContext_delay_54_payload_isFull <= fullRound_addContext_delay_53_payload_isFull;
    fullRound_addContext_delay_54_payload_fullRound <= fullRound_addContext_delay_53_payload_fullRound;
    fullRound_addContext_delay_54_payload_partialRound <= fullRound_addContext_delay_53_payload_partialRound;
    fullRound_addContext_delay_54_payload_stateSize <= fullRound_addContext_delay_53_payload_stateSize;
    fullRound_addContext_delay_54_payload_stateID <= fullRound_addContext_delay_53_payload_stateID;
    fullRound_addContext_delay_55_valid <= fullRound_addContext_delay_54_valid;
    fullRound_addContext_delay_55_payload_isFull <= fullRound_addContext_delay_54_payload_isFull;
    fullRound_addContext_delay_55_payload_fullRound <= fullRound_addContext_delay_54_payload_fullRound;
    fullRound_addContext_delay_55_payload_partialRound <= fullRound_addContext_delay_54_payload_partialRound;
    fullRound_addContext_delay_55_payload_stateSize <= fullRound_addContext_delay_54_payload_stateSize;
    fullRound_addContext_delay_55_payload_stateID <= fullRound_addContext_delay_54_payload_stateID;
    fullRound_addContext_delay_56_valid <= fullRound_addContext_delay_55_valid;
    fullRound_addContext_delay_56_payload_isFull <= fullRound_addContext_delay_55_payload_isFull;
    fullRound_addContext_delay_56_payload_fullRound <= fullRound_addContext_delay_55_payload_fullRound;
    fullRound_addContext_delay_56_payload_partialRound <= fullRound_addContext_delay_55_payload_partialRound;
    fullRound_addContext_delay_56_payload_stateSize <= fullRound_addContext_delay_55_payload_stateSize;
    fullRound_addContext_delay_56_payload_stateID <= fullRound_addContext_delay_55_payload_stateID;
    fullRound_addContext_delay_57_valid <= fullRound_addContext_delay_56_valid;
    fullRound_addContext_delay_57_payload_isFull <= fullRound_addContext_delay_56_payload_isFull;
    fullRound_addContext_delay_57_payload_fullRound <= fullRound_addContext_delay_56_payload_fullRound;
    fullRound_addContext_delay_57_payload_partialRound <= fullRound_addContext_delay_56_payload_partialRound;
    fullRound_addContext_delay_57_payload_stateSize <= fullRound_addContext_delay_56_payload_stateSize;
    fullRound_addContext_delay_57_payload_stateID <= fullRound_addContext_delay_56_payload_stateID;
    fullRound_addContext_delay_58_valid <= fullRound_addContext_delay_57_valid;
    fullRound_addContext_delay_58_payload_isFull <= fullRound_addContext_delay_57_payload_isFull;
    fullRound_addContext_delay_58_payload_fullRound <= fullRound_addContext_delay_57_payload_fullRound;
    fullRound_addContext_delay_58_payload_partialRound <= fullRound_addContext_delay_57_payload_partialRound;
    fullRound_addContext_delay_58_payload_stateSize <= fullRound_addContext_delay_57_payload_stateSize;
    fullRound_addContext_delay_58_payload_stateID <= fullRound_addContext_delay_57_payload_stateID;
    fullRound_addContext_delay_59_valid <= fullRound_addContext_delay_58_valid;
    fullRound_addContext_delay_59_payload_isFull <= fullRound_addContext_delay_58_payload_isFull;
    fullRound_addContext_delay_59_payload_fullRound <= fullRound_addContext_delay_58_payload_fullRound;
    fullRound_addContext_delay_59_payload_partialRound <= fullRound_addContext_delay_58_payload_partialRound;
    fullRound_addContext_delay_59_payload_stateSize <= fullRound_addContext_delay_58_payload_stateSize;
    fullRound_addContext_delay_59_payload_stateID <= fullRound_addContext_delay_58_payload_stateID;
    fullRound_addContext_delay_60_valid <= fullRound_addContext_delay_59_valid;
    fullRound_addContext_delay_60_payload_isFull <= fullRound_addContext_delay_59_payload_isFull;
    fullRound_addContext_delay_60_payload_fullRound <= fullRound_addContext_delay_59_payload_fullRound;
    fullRound_addContext_delay_60_payload_partialRound <= fullRound_addContext_delay_59_payload_partialRound;
    fullRound_addContext_delay_60_payload_stateSize <= fullRound_addContext_delay_59_payload_stateSize;
    fullRound_addContext_delay_60_payload_stateID <= fullRound_addContext_delay_59_payload_stateID;
    fullRound_addContext_delay_61_valid <= fullRound_addContext_delay_60_valid;
    fullRound_addContext_delay_61_payload_isFull <= fullRound_addContext_delay_60_payload_isFull;
    fullRound_addContext_delay_61_payload_fullRound <= fullRound_addContext_delay_60_payload_fullRound;
    fullRound_addContext_delay_61_payload_partialRound <= fullRound_addContext_delay_60_payload_partialRound;
    fullRound_addContext_delay_61_payload_stateSize <= fullRound_addContext_delay_60_payload_stateSize;
    fullRound_addContext_delay_61_payload_stateID <= fullRound_addContext_delay_60_payload_stateID;
    fullRound_addContext_delay_62_valid <= fullRound_addContext_delay_61_valid;
    fullRound_addContext_delay_62_payload_isFull <= fullRound_addContext_delay_61_payload_isFull;
    fullRound_addContext_delay_62_payload_fullRound <= fullRound_addContext_delay_61_payload_fullRound;
    fullRound_addContext_delay_62_payload_partialRound <= fullRound_addContext_delay_61_payload_partialRound;
    fullRound_addContext_delay_62_payload_stateSize <= fullRound_addContext_delay_61_payload_stateSize;
    fullRound_addContext_delay_62_payload_stateID <= fullRound_addContext_delay_61_payload_stateID;
    fullRound_addContext_delay_63_valid <= fullRound_addContext_delay_62_valid;
    fullRound_addContext_delay_63_payload_isFull <= fullRound_addContext_delay_62_payload_isFull;
    fullRound_addContext_delay_63_payload_fullRound <= fullRound_addContext_delay_62_payload_fullRound;
    fullRound_addContext_delay_63_payload_partialRound <= fullRound_addContext_delay_62_payload_partialRound;
    fullRound_addContext_delay_63_payload_stateSize <= fullRound_addContext_delay_62_payload_stateSize;
    fullRound_addContext_delay_63_payload_stateID <= fullRound_addContext_delay_62_payload_stateID;
    fullRound_addContextDelayed_valid <= fullRound_addContext_delay_63_valid;
    fullRound_addContextDelayed_payload_isFull <= fullRound_addContext_delay_63_payload_isFull;
    fullRound_addContextDelayed_payload_fullRound <= fullRound_addContext_delay_63_payload_fullRound;
    fullRound_addContextDelayed_payload_partialRound <= fullRound_addContext_delay_63_payload_partialRound;
    fullRound_addContextDelayed_payload_stateSize <= fullRound_addContext_delay_63_payload_stateSize;
    fullRound_addContextDelayed_payload_stateID <= fullRound_addContext_delay_63_payload_stateID;
    case(fullRound_deserialization_stateReg)
      fullRound_deserialization_enumDef_IDLE : begin
        if(fullRound_deserialization_adderTreeValid) begin
          fullRound_deserialization_tempOutput_isFull <= fullRound_addContextDelayed_payload_isFull;
          fullRound_deserialization_tempOutput_fullRound <= fullRound_addContextDelayed_payload_fullRound;
          fullRound_deserialization_tempOutput_partialRound <= fullRound_addContextDelayed_payload_partialRound;
          fullRound_deserialization_tempOutput_stateSize <= fullRound_addContextDelayed_payload_stateSize;
          fullRound_deserialization_tempOutput_stateID <= fullRound_addContextDelayed_payload_stateID;
        end
      end
      fullRound_deserialization_enumDef_BUSY : begin
      end
      fullRound_deserialization_enumDef_DONE : begin
        if(fullRound_deserialization_adderTreeValid) begin
          fullRound_deserialization_tempOutput_isFull <= fullRound_addContextDelayed_payload_isFull;
          fullRound_deserialization_tempOutput_fullRound <= fullRound_addContextDelayed_payload_fullRound;
          fullRound_deserialization_tempOutput_partialRound <= fullRound_addContextDelayed_payload_partialRound;
          fullRound_deserialization_tempOutput_stateSize <= fullRound_addContextDelayed_payload_stateSize;
          fullRound_deserialization_tempOutput_stateID <= fullRound_addContextDelayed_payload_stateID;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module MDSMatrixMultiplier (
  input               io_input_valid,
  input               io_input_payload_isFull,
  input      [2:0]    io_input_payload_fullRound,
  input      [5:0]    io_input_payload_partialRound,
  input      [3:0]    io_input_payload_stateIndex,
  input      [3:0]    io_input_payload_stateSize,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElements_0,
  input      [254:0]  io_input_payload_stateElements_1,
  input      [254:0]  io_input_payload_stateElements_2,
  input      [254:0]  io_input_payload_stateElements_3,
  input      [254:0]  io_input_payload_stateElements_4,
  input      [254:0]  io_input_payload_stateElements_5,
  input      [254:0]  io_input_payload_stateElements_6,
  input      [254:0]  io_input_payload_stateElements_7,
  input      [254:0]  io_input_payload_stateElements_8,
  input      [254:0]  io_input_payload_stateElements_9,
  input      [254:0]  io_input_payload_stateElements_10,
  input      [254:0]  io_input_payload_stateElement,
  output              io_output_valid,
  output              io_output_payload_isFull,
  output     [2:0]    io_output_payload_fullRound,
  output     [5:0]    io_output_payload_partialRound,
  output     [3:0]    io_output_payload_stateSize,
  output     [7:0]    io_output_payload_stateID,
  output     [254:0]  io_output_payload_stateElements_0,
  output     [254:0]  io_output_payload_stateElements_1,
  output     [254:0]  io_output_payload_stateElements_2,
  output     [254:0]  io_output_payload_stateElements_3,
  output     [254:0]  io_output_payload_stateElements_4,
  output     [254:0]  io_output_payload_stateElements_5,
  output     [254:0]  io_output_payload_stateElements_6,
  output     [254:0]  io_output_payload_stateElements_7,
  output     [254:0]  io_output_payload_stateElements_8,
  output     [254:0]  io_output_payload_stateElements_9,
  output     [254:0]  io_output_payload_stateElements_10,
  output     [254:0]  io_output_payload_stateElements_11,
  input               clk,
  input               resetn
);

  wire       [254:0]  constants_io_data_0;
  wire       [254:0]  constants_io_data_1;
  wire       [254:0]  constants_io_data_2;
  wire       [254:0]  constants_io_data_3;
  wire       [254:0]  constants_io_data_4;
  wire       [254:0]  constants_io_data_5;
  wire       [254:0]  constants_io_data_6;
  wire       [254:0]  constants_io_data_7;
  wire       [254:0]  constants_io_data_8;
  wire       [254:0]  constants_io_data_9;
  wire       [254:0]  constants_io_data_10;
  wire       [254:0]  constants_io_data_11;
  wire                montgomeryMultFlow_15_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_15_io_output_payload_res;
  wire                montgomeryMultFlow_16_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_16_io_output_payload_res;
  wire                montgomeryMultFlow_17_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_17_io_output_payload_res;
  wire                montgomeryMultFlow_18_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_18_io_output_payload_res;
  wire                montgomeryMultFlow_19_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_19_io_output_payload_res;
  wire                montgomeryMultFlow_20_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_20_io_output_payload_res;
  wire                montgomeryMultFlow_21_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_21_io_output_payload_res;
  wire                montgomeryMultFlow_22_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_22_io_output_payload_res;
  wire                montgomeryMultFlow_23_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_23_io_output_payload_res;
  wire                montgomeryMultFlow_24_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_24_io_output_payload_res;
  wire                montgomeryMultFlow_25_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_25_io_output_payload_res;
  wire                montgomeryMultFlow_26_io_output_valid;
  wire       [254:0]  montgomeryMultFlow_26_io_output_payload_res;
  wire       [254:0]  modAdderPiped_22_io_res;
  wire       [254:0]  modAdderPiped_23_io_res;
  wire       [254:0]  modAdderPiped_24_io_res;
  wire       [254:0]  modAdderPiped_25_io_res;
  wire       [254:0]  modAdderPiped_26_io_res;
  wire       [254:0]  modAdderPiped_27_io_res;
  wire       [254:0]  modAdderPiped_28_io_res;
  wire       [254:0]  modAdderPiped_29_io_res;
  wire       [254:0]  modAdderPiped_30_io_res;
  wire       [254:0]  modAdderPiped_31_io_res;
  wire       [254:0]  modAdderPiped_32_io_res;
  wire       [0:0]    _zz__zz_validDelayed;
  wire       [0:0]    _zz__zz_validDelayed_1;
  wire       [254:0]  _zz__zz_io_output_payload_stateElements_0;
  wire       [254:0]  _zz__zz_io_output_payload_stateElements_0_1;
  reg                 io_input_regNext_valid;
  reg                 io_input_regNext_payload_isFull;
  reg        [2:0]    io_input_regNext_payload_fullRound;
  reg        [5:0]    io_input_regNext_payload_partialRound;
  reg        [3:0]    io_input_regNext_payload_stateIndex;
  reg        [3:0]    io_input_regNext_payload_stateSize;
  reg        [7:0]    io_input_regNext_payload_stateID;
  reg        [254:0]  io_input_regNext_payload_stateElements_0;
  reg        [254:0]  io_input_regNext_payload_stateElements_1;
  reg        [254:0]  io_input_regNext_payload_stateElements_2;
  reg        [254:0]  io_input_regNext_payload_stateElements_3;
  reg        [254:0]  io_input_regNext_payload_stateElements_4;
  reg        [254:0]  io_input_regNext_payload_stateElements_5;
  reg        [254:0]  io_input_regNext_payload_stateElements_6;
  reg        [254:0]  io_input_regNext_payload_stateElements_7;
  reg        [254:0]  io_input_regNext_payload_stateElements_8;
  reg        [254:0]  io_input_regNext_payload_stateElements_9;
  reg        [254:0]  io_input_regNext_payload_stateElements_10;
  reg        [254:0]  io_input_regNext_payload_stateElement;
  reg                 io_input_regNext_regNext_valid;
  reg                 io_input_regNext_regNext_payload_isFull;
  reg        [2:0]    io_input_regNext_regNext_payload_fullRound;
  reg        [5:0]    io_input_regNext_regNext_payload_partialRound;
  reg        [3:0]    io_input_regNext_regNext_payload_stateIndex;
  reg        [3:0]    io_input_regNext_regNext_payload_stateSize;
  reg        [7:0]    io_input_regNext_regNext_payload_stateID;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_0;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_1;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_2;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_3;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_4;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_5;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_6;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_7;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_8;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_9;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElements_10;
  reg        [254:0]  io_input_regNext_regNext_payload_stateElement;
  reg                 io_input_regNext_regNext_regNext_valid;
  reg                 io_input_regNext_regNext_regNext_payload_isFull;
  reg        [2:0]    io_input_regNext_regNext_regNext_payload_fullRound;
  reg        [5:0]    io_input_regNext_regNext_regNext_payload_partialRound;
  reg        [3:0]    io_input_regNext_regNext_regNext_payload_stateIndex;
  reg        [3:0]    io_input_regNext_regNext_regNext_payload_stateSize;
  reg        [7:0]    io_input_regNext_regNext_regNext_payload_stateID;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_0;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_1;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_2;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_3;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_4;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_5;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_6;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_7;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_8;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_9;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElements_10;
  reg        [254:0]  io_input_regNext_regNext_regNext_payload_stateElement;
  reg                 io_input_regNext_regNext_regNext_regNext_valid;
  reg                 io_input_regNext_regNext_regNext_regNext_payload_isFull;
  reg        [2:0]    io_input_regNext_regNext_regNext_regNext_payload_fullRound;
  reg        [5:0]    io_input_regNext_regNext_regNext_regNext_payload_partialRound;
  reg        [3:0]    io_input_regNext_regNext_regNext_regNext_payload_stateIndex;
  reg        [3:0]    io_input_regNext_regNext_regNext_regNext_payload_stateSize;
  reg        [7:0]    io_input_regNext_regNext_regNext_regNext_payload_stateID;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_0;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_1;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_2;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_3;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_4;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_5;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_6;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_7;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_8;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_9;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElements_10;
  reg        [254:0]  io_input_regNext_regNext_regNext_regNext_payload_stateElement;
  reg                 inputDelayed_valid;
  reg                 inputDelayed_payload_isFull;
  reg        [2:0]    inputDelayed_payload_fullRound;
  reg        [5:0]    inputDelayed_payload_partialRound;
  reg        [3:0]    inputDelayed_payload_stateIndex;
  reg        [3:0]    inputDelayed_payload_stateSize;
  reg        [7:0]    inputDelayed_payload_stateID;
  reg        [254:0]  inputDelayed_payload_stateElements_0;
  reg        [254:0]  inputDelayed_payload_stateElements_1;
  reg        [254:0]  inputDelayed_payload_stateElements_2;
  reg        [254:0]  inputDelayed_payload_stateElements_3;
  reg        [254:0]  inputDelayed_payload_stateElements_4;
  reg        [254:0]  inputDelayed_payload_stateElements_5;
  reg        [254:0]  inputDelayed_payload_stateElements_6;
  reg        [254:0]  inputDelayed_payload_stateElements_7;
  reg        [254:0]  inputDelayed_payload_stateElements_8;
  reg        [254:0]  inputDelayed_payload_stateElements_9;
  reg        [254:0]  inputDelayed_payload_stateElements_10;
  reg        [254:0]  inputDelayed_payload_stateElement;
  wire                mulInputs_0_valid;
  wire       [254:0]  mulInputs_0_payload_op1;
  wire       [254:0]  mulInputs_0_payload_op2;
  wire                mulInputs_1_valid;
  reg        [254:0]  mulInputs_1_payload_op1;
  wire       [254:0]  mulInputs_1_payload_op2;
  wire                mulInputs_2_valid;
  reg        [254:0]  mulInputs_2_payload_op1;
  wire       [254:0]  mulInputs_2_payload_op2;
  wire                mulInputs_3_valid;
  reg        [254:0]  mulInputs_3_payload_op1;
  wire       [254:0]  mulInputs_3_payload_op2;
  wire                mulInputs_4_valid;
  reg        [254:0]  mulInputs_4_payload_op1;
  wire       [254:0]  mulInputs_4_payload_op2;
  wire                mulInputs_5_valid;
  reg        [254:0]  mulInputs_5_payload_op1;
  wire       [254:0]  mulInputs_5_payload_op2;
  wire                mulInputs_6_valid;
  reg        [254:0]  mulInputs_6_payload_op1;
  wire       [254:0]  mulInputs_6_payload_op2;
  wire                mulInputs_7_valid;
  reg        [254:0]  mulInputs_7_payload_op1;
  wire       [254:0]  mulInputs_7_payload_op2;
  wire                mulInputs_8_valid;
  reg        [254:0]  mulInputs_8_payload_op1;
  wire       [254:0]  mulInputs_8_payload_op2;
  wire                mulInputs_9_valid;
  reg        [254:0]  mulInputs_9_payload_op1;
  wire       [254:0]  mulInputs_9_payload_op2;
  wire                mulInputs_10_valid;
  reg        [254:0]  mulInputs_10_payload_op1;
  wire       [254:0]  mulInputs_10_payload_op2;
  wire                mulInputs_11_valid;
  reg        [254:0]  mulInputs_11_payload_op1;
  wire       [254:0]  mulInputs_11_payload_op2;
  wire                when_MDSMatrixMultiplier_l73;
  wire                when_MDSMatrixMultiplier_l74;
  wire                when_MDSMatrixMultiplier_l76;
  wire                when_MDSMatrixMultiplier_l78;
  reg                 mulInputsTemp_0_valid;
  reg        [254:0]  mulInputsTemp_0_payload_op1;
  reg        [254:0]  mulInputsTemp_0_payload_op2;
  reg                 mulInputsTemp_1_valid;
  reg        [254:0]  mulInputsTemp_1_payload_op1;
  reg        [254:0]  mulInputsTemp_1_payload_op2;
  reg                 mulInputsTemp_2_valid;
  reg        [254:0]  mulInputsTemp_2_payload_op1;
  reg        [254:0]  mulInputsTemp_2_payload_op2;
  reg                 mulInputsTemp_3_valid;
  reg        [254:0]  mulInputsTemp_3_payload_op1;
  reg        [254:0]  mulInputsTemp_3_payload_op2;
  reg                 mulInputsTemp_4_valid;
  reg        [254:0]  mulInputsTemp_4_payload_op1;
  reg        [254:0]  mulInputsTemp_4_payload_op2;
  reg                 mulInputsTemp_5_valid;
  reg        [254:0]  mulInputsTemp_5_payload_op1;
  reg        [254:0]  mulInputsTemp_5_payload_op2;
  reg                 mulInputsTemp_6_valid;
  reg        [254:0]  mulInputsTemp_6_payload_op1;
  reg        [254:0]  mulInputsTemp_6_payload_op2;
  reg                 mulInputsTemp_7_valid;
  reg        [254:0]  mulInputsTemp_7_payload_op1;
  reg        [254:0]  mulInputsTemp_7_payload_op2;
  reg                 mulInputsTemp_8_valid;
  reg        [254:0]  mulInputsTemp_8_payload_op1;
  reg        [254:0]  mulInputsTemp_8_payload_op2;
  reg                 mulInputsTemp_9_valid;
  reg        [254:0]  mulInputsTemp_9_payload_op1;
  reg        [254:0]  mulInputsTemp_9_payload_op2;
  reg                 mulInputsTemp_10_valid;
  reg        [254:0]  mulInputsTemp_10_payload_op1;
  reg        [254:0]  mulInputsTemp_10_payload_op2;
  reg                 mulInputsTemp_11_valid;
  reg        [254:0]  mulInputsTemp_11_payload_op1;
  reg        [254:0]  mulInputsTemp_11_payload_op2;
  wire                mulContext_isFull;
  wire       [2:0]    mulContext_fullRound;
  wire       [5:0]    mulContext_partialRound;
  wire       [3:0]    mulContext_stateSize;
  wire       [7:0]    mulContext_stateID;
  reg        [254:0]  mulContext_stateElements_0;
  reg        [254:0]  mulContext_stateElements_1;
  reg        [254:0]  mulContext_stateElements_2;
  reg        [254:0]  mulContext_stateElements_3;
  reg        [254:0]  mulContext_stateElements_4;
  reg        [254:0]  mulContext_stateElements_5;
  reg        [254:0]  mulContext_stateElements_6;
  reg        [254:0]  mulContext_stateElements_7;
  reg        [254:0]  mulContext_stateElements_8;
  reg        [254:0]  mulContext_stateElements_9;
  reg        [254:0]  mulContext_stateElements_10;
  wire                when_MDSMatrixMultiplier_l94;
  wire       [2804:0] _zz_mulContext_stateElements_0;
  reg                 mulContext_delay_1_isFull;
  reg        [2:0]    mulContext_delay_1_fullRound;
  reg        [5:0]    mulContext_delay_1_partialRound;
  reg        [3:0]    mulContext_delay_1_stateSize;
  reg        [7:0]    mulContext_delay_1_stateID;
  reg        [254:0]  mulContext_delay_1_stateElements_0;
  reg        [254:0]  mulContext_delay_1_stateElements_1;
  reg        [254:0]  mulContext_delay_1_stateElements_2;
  reg        [254:0]  mulContext_delay_1_stateElements_3;
  reg        [254:0]  mulContext_delay_1_stateElements_4;
  reg        [254:0]  mulContext_delay_1_stateElements_5;
  reg        [254:0]  mulContext_delay_1_stateElements_6;
  reg        [254:0]  mulContext_delay_1_stateElements_7;
  reg        [254:0]  mulContext_delay_1_stateElements_8;
  reg        [254:0]  mulContext_delay_1_stateElements_9;
  reg        [254:0]  mulContext_delay_1_stateElements_10;
  reg                 mulContext_delay_2_isFull;
  reg        [2:0]    mulContext_delay_2_fullRound;
  reg        [5:0]    mulContext_delay_2_partialRound;
  reg        [3:0]    mulContext_delay_2_stateSize;
  reg        [7:0]    mulContext_delay_2_stateID;
  reg        [254:0]  mulContext_delay_2_stateElements_0;
  reg        [254:0]  mulContext_delay_2_stateElements_1;
  reg        [254:0]  mulContext_delay_2_stateElements_2;
  reg        [254:0]  mulContext_delay_2_stateElements_3;
  reg        [254:0]  mulContext_delay_2_stateElements_4;
  reg        [254:0]  mulContext_delay_2_stateElements_5;
  reg        [254:0]  mulContext_delay_2_stateElements_6;
  reg        [254:0]  mulContext_delay_2_stateElements_7;
  reg        [254:0]  mulContext_delay_2_stateElements_8;
  reg        [254:0]  mulContext_delay_2_stateElements_9;
  reg        [254:0]  mulContext_delay_2_stateElements_10;
  reg                 mulContext_delay_3_isFull;
  reg        [2:0]    mulContext_delay_3_fullRound;
  reg        [5:0]    mulContext_delay_3_partialRound;
  reg        [3:0]    mulContext_delay_3_stateSize;
  reg        [7:0]    mulContext_delay_3_stateID;
  reg        [254:0]  mulContext_delay_3_stateElements_0;
  reg        [254:0]  mulContext_delay_3_stateElements_1;
  reg        [254:0]  mulContext_delay_3_stateElements_2;
  reg        [254:0]  mulContext_delay_3_stateElements_3;
  reg        [254:0]  mulContext_delay_3_stateElements_4;
  reg        [254:0]  mulContext_delay_3_stateElements_5;
  reg        [254:0]  mulContext_delay_3_stateElements_6;
  reg        [254:0]  mulContext_delay_3_stateElements_7;
  reg        [254:0]  mulContext_delay_3_stateElements_8;
  reg        [254:0]  mulContext_delay_3_stateElements_9;
  reg        [254:0]  mulContext_delay_3_stateElements_10;
  reg                 mulContext_delay_4_isFull;
  reg        [2:0]    mulContext_delay_4_fullRound;
  reg        [5:0]    mulContext_delay_4_partialRound;
  reg        [3:0]    mulContext_delay_4_stateSize;
  reg        [7:0]    mulContext_delay_4_stateID;
  reg        [254:0]  mulContext_delay_4_stateElements_0;
  reg        [254:0]  mulContext_delay_4_stateElements_1;
  reg        [254:0]  mulContext_delay_4_stateElements_2;
  reg        [254:0]  mulContext_delay_4_stateElements_3;
  reg        [254:0]  mulContext_delay_4_stateElements_4;
  reg        [254:0]  mulContext_delay_4_stateElements_5;
  reg        [254:0]  mulContext_delay_4_stateElements_6;
  reg        [254:0]  mulContext_delay_4_stateElements_7;
  reg        [254:0]  mulContext_delay_4_stateElements_8;
  reg        [254:0]  mulContext_delay_4_stateElements_9;
  reg        [254:0]  mulContext_delay_4_stateElements_10;
  reg                 mulContext_delay_5_isFull;
  reg        [2:0]    mulContext_delay_5_fullRound;
  reg        [5:0]    mulContext_delay_5_partialRound;
  reg        [3:0]    mulContext_delay_5_stateSize;
  reg        [7:0]    mulContext_delay_5_stateID;
  reg        [254:0]  mulContext_delay_5_stateElements_0;
  reg        [254:0]  mulContext_delay_5_stateElements_1;
  reg        [254:0]  mulContext_delay_5_stateElements_2;
  reg        [254:0]  mulContext_delay_5_stateElements_3;
  reg        [254:0]  mulContext_delay_5_stateElements_4;
  reg        [254:0]  mulContext_delay_5_stateElements_5;
  reg        [254:0]  mulContext_delay_5_stateElements_6;
  reg        [254:0]  mulContext_delay_5_stateElements_7;
  reg        [254:0]  mulContext_delay_5_stateElements_8;
  reg        [254:0]  mulContext_delay_5_stateElements_9;
  reg        [254:0]  mulContext_delay_5_stateElements_10;
  reg                 mulContext_delay_6_isFull;
  reg        [2:0]    mulContext_delay_6_fullRound;
  reg        [5:0]    mulContext_delay_6_partialRound;
  reg        [3:0]    mulContext_delay_6_stateSize;
  reg        [7:0]    mulContext_delay_6_stateID;
  reg        [254:0]  mulContext_delay_6_stateElements_0;
  reg        [254:0]  mulContext_delay_6_stateElements_1;
  reg        [254:0]  mulContext_delay_6_stateElements_2;
  reg        [254:0]  mulContext_delay_6_stateElements_3;
  reg        [254:0]  mulContext_delay_6_stateElements_4;
  reg        [254:0]  mulContext_delay_6_stateElements_5;
  reg        [254:0]  mulContext_delay_6_stateElements_6;
  reg        [254:0]  mulContext_delay_6_stateElements_7;
  reg        [254:0]  mulContext_delay_6_stateElements_8;
  reg        [254:0]  mulContext_delay_6_stateElements_9;
  reg        [254:0]  mulContext_delay_6_stateElements_10;
  reg                 mulContext_delay_7_isFull;
  reg        [2:0]    mulContext_delay_7_fullRound;
  reg        [5:0]    mulContext_delay_7_partialRound;
  reg        [3:0]    mulContext_delay_7_stateSize;
  reg        [7:0]    mulContext_delay_7_stateID;
  reg        [254:0]  mulContext_delay_7_stateElements_0;
  reg        [254:0]  mulContext_delay_7_stateElements_1;
  reg        [254:0]  mulContext_delay_7_stateElements_2;
  reg        [254:0]  mulContext_delay_7_stateElements_3;
  reg        [254:0]  mulContext_delay_7_stateElements_4;
  reg        [254:0]  mulContext_delay_7_stateElements_5;
  reg        [254:0]  mulContext_delay_7_stateElements_6;
  reg        [254:0]  mulContext_delay_7_stateElements_7;
  reg        [254:0]  mulContext_delay_7_stateElements_8;
  reg        [254:0]  mulContext_delay_7_stateElements_9;
  reg        [254:0]  mulContext_delay_7_stateElements_10;
  reg                 mulContext_delay_8_isFull;
  reg        [2:0]    mulContext_delay_8_fullRound;
  reg        [5:0]    mulContext_delay_8_partialRound;
  reg        [3:0]    mulContext_delay_8_stateSize;
  reg        [7:0]    mulContext_delay_8_stateID;
  reg        [254:0]  mulContext_delay_8_stateElements_0;
  reg        [254:0]  mulContext_delay_8_stateElements_1;
  reg        [254:0]  mulContext_delay_8_stateElements_2;
  reg        [254:0]  mulContext_delay_8_stateElements_3;
  reg        [254:0]  mulContext_delay_8_stateElements_4;
  reg        [254:0]  mulContext_delay_8_stateElements_5;
  reg        [254:0]  mulContext_delay_8_stateElements_6;
  reg        [254:0]  mulContext_delay_8_stateElements_7;
  reg        [254:0]  mulContext_delay_8_stateElements_8;
  reg        [254:0]  mulContext_delay_8_stateElements_9;
  reg        [254:0]  mulContext_delay_8_stateElements_10;
  reg                 mulContext_delay_9_isFull;
  reg        [2:0]    mulContext_delay_9_fullRound;
  reg        [5:0]    mulContext_delay_9_partialRound;
  reg        [3:0]    mulContext_delay_9_stateSize;
  reg        [7:0]    mulContext_delay_9_stateID;
  reg        [254:0]  mulContext_delay_9_stateElements_0;
  reg        [254:0]  mulContext_delay_9_stateElements_1;
  reg        [254:0]  mulContext_delay_9_stateElements_2;
  reg        [254:0]  mulContext_delay_9_stateElements_3;
  reg        [254:0]  mulContext_delay_9_stateElements_4;
  reg        [254:0]  mulContext_delay_9_stateElements_5;
  reg        [254:0]  mulContext_delay_9_stateElements_6;
  reg        [254:0]  mulContext_delay_9_stateElements_7;
  reg        [254:0]  mulContext_delay_9_stateElements_8;
  reg        [254:0]  mulContext_delay_9_stateElements_9;
  reg        [254:0]  mulContext_delay_9_stateElements_10;
  reg                 mulContext_delay_10_isFull;
  reg        [2:0]    mulContext_delay_10_fullRound;
  reg        [5:0]    mulContext_delay_10_partialRound;
  reg        [3:0]    mulContext_delay_10_stateSize;
  reg        [7:0]    mulContext_delay_10_stateID;
  reg        [254:0]  mulContext_delay_10_stateElements_0;
  reg        [254:0]  mulContext_delay_10_stateElements_1;
  reg        [254:0]  mulContext_delay_10_stateElements_2;
  reg        [254:0]  mulContext_delay_10_stateElements_3;
  reg        [254:0]  mulContext_delay_10_stateElements_4;
  reg        [254:0]  mulContext_delay_10_stateElements_5;
  reg        [254:0]  mulContext_delay_10_stateElements_6;
  reg        [254:0]  mulContext_delay_10_stateElements_7;
  reg        [254:0]  mulContext_delay_10_stateElements_8;
  reg        [254:0]  mulContext_delay_10_stateElements_9;
  reg        [254:0]  mulContext_delay_10_stateElements_10;
  reg                 mulContext_delay_11_isFull;
  reg        [2:0]    mulContext_delay_11_fullRound;
  reg        [5:0]    mulContext_delay_11_partialRound;
  reg        [3:0]    mulContext_delay_11_stateSize;
  reg        [7:0]    mulContext_delay_11_stateID;
  reg        [254:0]  mulContext_delay_11_stateElements_0;
  reg        [254:0]  mulContext_delay_11_stateElements_1;
  reg        [254:0]  mulContext_delay_11_stateElements_2;
  reg        [254:0]  mulContext_delay_11_stateElements_3;
  reg        [254:0]  mulContext_delay_11_stateElements_4;
  reg        [254:0]  mulContext_delay_11_stateElements_5;
  reg        [254:0]  mulContext_delay_11_stateElements_6;
  reg        [254:0]  mulContext_delay_11_stateElements_7;
  reg        [254:0]  mulContext_delay_11_stateElements_8;
  reg        [254:0]  mulContext_delay_11_stateElements_9;
  reg        [254:0]  mulContext_delay_11_stateElements_10;
  reg                 mulContext_delay_12_isFull;
  reg        [2:0]    mulContext_delay_12_fullRound;
  reg        [5:0]    mulContext_delay_12_partialRound;
  reg        [3:0]    mulContext_delay_12_stateSize;
  reg        [7:0]    mulContext_delay_12_stateID;
  reg        [254:0]  mulContext_delay_12_stateElements_0;
  reg        [254:0]  mulContext_delay_12_stateElements_1;
  reg        [254:0]  mulContext_delay_12_stateElements_2;
  reg        [254:0]  mulContext_delay_12_stateElements_3;
  reg        [254:0]  mulContext_delay_12_stateElements_4;
  reg        [254:0]  mulContext_delay_12_stateElements_5;
  reg        [254:0]  mulContext_delay_12_stateElements_6;
  reg        [254:0]  mulContext_delay_12_stateElements_7;
  reg        [254:0]  mulContext_delay_12_stateElements_8;
  reg        [254:0]  mulContext_delay_12_stateElements_9;
  reg        [254:0]  mulContext_delay_12_stateElements_10;
  reg                 mulContext_delay_13_isFull;
  reg        [2:0]    mulContext_delay_13_fullRound;
  reg        [5:0]    mulContext_delay_13_partialRound;
  reg        [3:0]    mulContext_delay_13_stateSize;
  reg        [7:0]    mulContext_delay_13_stateID;
  reg        [254:0]  mulContext_delay_13_stateElements_0;
  reg        [254:0]  mulContext_delay_13_stateElements_1;
  reg        [254:0]  mulContext_delay_13_stateElements_2;
  reg        [254:0]  mulContext_delay_13_stateElements_3;
  reg        [254:0]  mulContext_delay_13_stateElements_4;
  reg        [254:0]  mulContext_delay_13_stateElements_5;
  reg        [254:0]  mulContext_delay_13_stateElements_6;
  reg        [254:0]  mulContext_delay_13_stateElements_7;
  reg        [254:0]  mulContext_delay_13_stateElements_8;
  reg        [254:0]  mulContext_delay_13_stateElements_9;
  reg        [254:0]  mulContext_delay_13_stateElements_10;
  reg                 mulContext_delay_14_isFull;
  reg        [2:0]    mulContext_delay_14_fullRound;
  reg        [5:0]    mulContext_delay_14_partialRound;
  reg        [3:0]    mulContext_delay_14_stateSize;
  reg        [7:0]    mulContext_delay_14_stateID;
  reg        [254:0]  mulContext_delay_14_stateElements_0;
  reg        [254:0]  mulContext_delay_14_stateElements_1;
  reg        [254:0]  mulContext_delay_14_stateElements_2;
  reg        [254:0]  mulContext_delay_14_stateElements_3;
  reg        [254:0]  mulContext_delay_14_stateElements_4;
  reg        [254:0]  mulContext_delay_14_stateElements_5;
  reg        [254:0]  mulContext_delay_14_stateElements_6;
  reg        [254:0]  mulContext_delay_14_stateElements_7;
  reg        [254:0]  mulContext_delay_14_stateElements_8;
  reg        [254:0]  mulContext_delay_14_stateElements_9;
  reg        [254:0]  mulContext_delay_14_stateElements_10;
  reg                 mulContext_delay_15_isFull;
  reg        [2:0]    mulContext_delay_15_fullRound;
  reg        [5:0]    mulContext_delay_15_partialRound;
  reg        [3:0]    mulContext_delay_15_stateSize;
  reg        [7:0]    mulContext_delay_15_stateID;
  reg        [254:0]  mulContext_delay_15_stateElements_0;
  reg        [254:0]  mulContext_delay_15_stateElements_1;
  reg        [254:0]  mulContext_delay_15_stateElements_2;
  reg        [254:0]  mulContext_delay_15_stateElements_3;
  reg        [254:0]  mulContext_delay_15_stateElements_4;
  reg        [254:0]  mulContext_delay_15_stateElements_5;
  reg        [254:0]  mulContext_delay_15_stateElements_6;
  reg        [254:0]  mulContext_delay_15_stateElements_7;
  reg        [254:0]  mulContext_delay_15_stateElements_8;
  reg        [254:0]  mulContext_delay_15_stateElements_9;
  reg        [254:0]  mulContext_delay_15_stateElements_10;
  reg                 mulContext_delay_16_isFull;
  reg        [2:0]    mulContext_delay_16_fullRound;
  reg        [5:0]    mulContext_delay_16_partialRound;
  reg        [3:0]    mulContext_delay_16_stateSize;
  reg        [7:0]    mulContext_delay_16_stateID;
  reg        [254:0]  mulContext_delay_16_stateElements_0;
  reg        [254:0]  mulContext_delay_16_stateElements_1;
  reg        [254:0]  mulContext_delay_16_stateElements_2;
  reg        [254:0]  mulContext_delay_16_stateElements_3;
  reg        [254:0]  mulContext_delay_16_stateElements_4;
  reg        [254:0]  mulContext_delay_16_stateElements_5;
  reg        [254:0]  mulContext_delay_16_stateElements_6;
  reg        [254:0]  mulContext_delay_16_stateElements_7;
  reg        [254:0]  mulContext_delay_16_stateElements_8;
  reg        [254:0]  mulContext_delay_16_stateElements_9;
  reg        [254:0]  mulContext_delay_16_stateElements_10;
  reg                 mulContext_delay_17_isFull;
  reg        [2:0]    mulContext_delay_17_fullRound;
  reg        [5:0]    mulContext_delay_17_partialRound;
  reg        [3:0]    mulContext_delay_17_stateSize;
  reg        [7:0]    mulContext_delay_17_stateID;
  reg        [254:0]  mulContext_delay_17_stateElements_0;
  reg        [254:0]  mulContext_delay_17_stateElements_1;
  reg        [254:0]  mulContext_delay_17_stateElements_2;
  reg        [254:0]  mulContext_delay_17_stateElements_3;
  reg        [254:0]  mulContext_delay_17_stateElements_4;
  reg        [254:0]  mulContext_delay_17_stateElements_5;
  reg        [254:0]  mulContext_delay_17_stateElements_6;
  reg        [254:0]  mulContext_delay_17_stateElements_7;
  reg        [254:0]  mulContext_delay_17_stateElements_8;
  reg        [254:0]  mulContext_delay_17_stateElements_9;
  reg        [254:0]  mulContext_delay_17_stateElements_10;
  reg                 mulContext_delay_18_isFull;
  reg        [2:0]    mulContext_delay_18_fullRound;
  reg        [5:0]    mulContext_delay_18_partialRound;
  reg        [3:0]    mulContext_delay_18_stateSize;
  reg        [7:0]    mulContext_delay_18_stateID;
  reg        [254:0]  mulContext_delay_18_stateElements_0;
  reg        [254:0]  mulContext_delay_18_stateElements_1;
  reg        [254:0]  mulContext_delay_18_stateElements_2;
  reg        [254:0]  mulContext_delay_18_stateElements_3;
  reg        [254:0]  mulContext_delay_18_stateElements_4;
  reg        [254:0]  mulContext_delay_18_stateElements_5;
  reg        [254:0]  mulContext_delay_18_stateElements_6;
  reg        [254:0]  mulContext_delay_18_stateElements_7;
  reg        [254:0]  mulContext_delay_18_stateElements_8;
  reg        [254:0]  mulContext_delay_18_stateElements_9;
  reg        [254:0]  mulContext_delay_18_stateElements_10;
  reg                 mulContext_delay_19_isFull;
  reg        [2:0]    mulContext_delay_19_fullRound;
  reg        [5:0]    mulContext_delay_19_partialRound;
  reg        [3:0]    mulContext_delay_19_stateSize;
  reg        [7:0]    mulContext_delay_19_stateID;
  reg        [254:0]  mulContext_delay_19_stateElements_0;
  reg        [254:0]  mulContext_delay_19_stateElements_1;
  reg        [254:0]  mulContext_delay_19_stateElements_2;
  reg        [254:0]  mulContext_delay_19_stateElements_3;
  reg        [254:0]  mulContext_delay_19_stateElements_4;
  reg        [254:0]  mulContext_delay_19_stateElements_5;
  reg        [254:0]  mulContext_delay_19_stateElements_6;
  reg        [254:0]  mulContext_delay_19_stateElements_7;
  reg        [254:0]  mulContext_delay_19_stateElements_8;
  reg        [254:0]  mulContext_delay_19_stateElements_9;
  reg        [254:0]  mulContext_delay_19_stateElements_10;
  reg                 mulContext_delay_20_isFull;
  reg        [2:0]    mulContext_delay_20_fullRound;
  reg        [5:0]    mulContext_delay_20_partialRound;
  reg        [3:0]    mulContext_delay_20_stateSize;
  reg        [7:0]    mulContext_delay_20_stateID;
  reg        [254:0]  mulContext_delay_20_stateElements_0;
  reg        [254:0]  mulContext_delay_20_stateElements_1;
  reg        [254:0]  mulContext_delay_20_stateElements_2;
  reg        [254:0]  mulContext_delay_20_stateElements_3;
  reg        [254:0]  mulContext_delay_20_stateElements_4;
  reg        [254:0]  mulContext_delay_20_stateElements_5;
  reg        [254:0]  mulContext_delay_20_stateElements_6;
  reg        [254:0]  mulContext_delay_20_stateElements_7;
  reg        [254:0]  mulContext_delay_20_stateElements_8;
  reg        [254:0]  mulContext_delay_20_stateElements_9;
  reg        [254:0]  mulContext_delay_20_stateElements_10;
  reg                 mulContext_delay_21_isFull;
  reg        [2:0]    mulContext_delay_21_fullRound;
  reg        [5:0]    mulContext_delay_21_partialRound;
  reg        [3:0]    mulContext_delay_21_stateSize;
  reg        [7:0]    mulContext_delay_21_stateID;
  reg        [254:0]  mulContext_delay_21_stateElements_0;
  reg        [254:0]  mulContext_delay_21_stateElements_1;
  reg        [254:0]  mulContext_delay_21_stateElements_2;
  reg        [254:0]  mulContext_delay_21_stateElements_3;
  reg        [254:0]  mulContext_delay_21_stateElements_4;
  reg        [254:0]  mulContext_delay_21_stateElements_5;
  reg        [254:0]  mulContext_delay_21_stateElements_6;
  reg        [254:0]  mulContext_delay_21_stateElements_7;
  reg        [254:0]  mulContext_delay_21_stateElements_8;
  reg        [254:0]  mulContext_delay_21_stateElements_9;
  reg        [254:0]  mulContext_delay_21_stateElements_10;
  reg                 mulContext_delay_22_isFull;
  reg        [2:0]    mulContext_delay_22_fullRound;
  reg        [5:0]    mulContext_delay_22_partialRound;
  reg        [3:0]    mulContext_delay_22_stateSize;
  reg        [7:0]    mulContext_delay_22_stateID;
  reg        [254:0]  mulContext_delay_22_stateElements_0;
  reg        [254:0]  mulContext_delay_22_stateElements_1;
  reg        [254:0]  mulContext_delay_22_stateElements_2;
  reg        [254:0]  mulContext_delay_22_stateElements_3;
  reg        [254:0]  mulContext_delay_22_stateElements_4;
  reg        [254:0]  mulContext_delay_22_stateElements_5;
  reg        [254:0]  mulContext_delay_22_stateElements_6;
  reg        [254:0]  mulContext_delay_22_stateElements_7;
  reg        [254:0]  mulContext_delay_22_stateElements_8;
  reg        [254:0]  mulContext_delay_22_stateElements_9;
  reg        [254:0]  mulContext_delay_22_stateElements_10;
  reg                 mulContext_delay_23_isFull;
  reg        [2:0]    mulContext_delay_23_fullRound;
  reg        [5:0]    mulContext_delay_23_partialRound;
  reg        [3:0]    mulContext_delay_23_stateSize;
  reg        [7:0]    mulContext_delay_23_stateID;
  reg        [254:0]  mulContext_delay_23_stateElements_0;
  reg        [254:0]  mulContext_delay_23_stateElements_1;
  reg        [254:0]  mulContext_delay_23_stateElements_2;
  reg        [254:0]  mulContext_delay_23_stateElements_3;
  reg        [254:0]  mulContext_delay_23_stateElements_4;
  reg        [254:0]  mulContext_delay_23_stateElements_5;
  reg        [254:0]  mulContext_delay_23_stateElements_6;
  reg        [254:0]  mulContext_delay_23_stateElements_7;
  reg        [254:0]  mulContext_delay_23_stateElements_8;
  reg        [254:0]  mulContext_delay_23_stateElements_9;
  reg        [254:0]  mulContext_delay_23_stateElements_10;
  reg                 mulContext_delay_24_isFull;
  reg        [2:0]    mulContext_delay_24_fullRound;
  reg        [5:0]    mulContext_delay_24_partialRound;
  reg        [3:0]    mulContext_delay_24_stateSize;
  reg        [7:0]    mulContext_delay_24_stateID;
  reg        [254:0]  mulContext_delay_24_stateElements_0;
  reg        [254:0]  mulContext_delay_24_stateElements_1;
  reg        [254:0]  mulContext_delay_24_stateElements_2;
  reg        [254:0]  mulContext_delay_24_stateElements_3;
  reg        [254:0]  mulContext_delay_24_stateElements_4;
  reg        [254:0]  mulContext_delay_24_stateElements_5;
  reg        [254:0]  mulContext_delay_24_stateElements_6;
  reg        [254:0]  mulContext_delay_24_stateElements_7;
  reg        [254:0]  mulContext_delay_24_stateElements_8;
  reg        [254:0]  mulContext_delay_24_stateElements_9;
  reg        [254:0]  mulContext_delay_24_stateElements_10;
  reg                 mulContext_delay_25_isFull;
  reg        [2:0]    mulContext_delay_25_fullRound;
  reg        [5:0]    mulContext_delay_25_partialRound;
  reg        [3:0]    mulContext_delay_25_stateSize;
  reg        [7:0]    mulContext_delay_25_stateID;
  reg        [254:0]  mulContext_delay_25_stateElements_0;
  reg        [254:0]  mulContext_delay_25_stateElements_1;
  reg        [254:0]  mulContext_delay_25_stateElements_2;
  reg        [254:0]  mulContext_delay_25_stateElements_3;
  reg        [254:0]  mulContext_delay_25_stateElements_4;
  reg        [254:0]  mulContext_delay_25_stateElements_5;
  reg        [254:0]  mulContext_delay_25_stateElements_6;
  reg        [254:0]  mulContext_delay_25_stateElements_7;
  reg        [254:0]  mulContext_delay_25_stateElements_8;
  reg        [254:0]  mulContext_delay_25_stateElements_9;
  reg        [254:0]  mulContext_delay_25_stateElements_10;
  reg                 mulContext_delay_26_isFull;
  reg        [2:0]    mulContext_delay_26_fullRound;
  reg        [5:0]    mulContext_delay_26_partialRound;
  reg        [3:0]    mulContext_delay_26_stateSize;
  reg        [7:0]    mulContext_delay_26_stateID;
  reg        [254:0]  mulContext_delay_26_stateElements_0;
  reg        [254:0]  mulContext_delay_26_stateElements_1;
  reg        [254:0]  mulContext_delay_26_stateElements_2;
  reg        [254:0]  mulContext_delay_26_stateElements_3;
  reg        [254:0]  mulContext_delay_26_stateElements_4;
  reg        [254:0]  mulContext_delay_26_stateElements_5;
  reg        [254:0]  mulContext_delay_26_stateElements_6;
  reg        [254:0]  mulContext_delay_26_stateElements_7;
  reg        [254:0]  mulContext_delay_26_stateElements_8;
  reg        [254:0]  mulContext_delay_26_stateElements_9;
  reg        [254:0]  mulContext_delay_26_stateElements_10;
  reg                 mulContext_delay_27_isFull;
  reg        [2:0]    mulContext_delay_27_fullRound;
  reg        [5:0]    mulContext_delay_27_partialRound;
  reg        [3:0]    mulContext_delay_27_stateSize;
  reg        [7:0]    mulContext_delay_27_stateID;
  reg        [254:0]  mulContext_delay_27_stateElements_0;
  reg        [254:0]  mulContext_delay_27_stateElements_1;
  reg        [254:0]  mulContext_delay_27_stateElements_2;
  reg        [254:0]  mulContext_delay_27_stateElements_3;
  reg        [254:0]  mulContext_delay_27_stateElements_4;
  reg        [254:0]  mulContext_delay_27_stateElements_5;
  reg        [254:0]  mulContext_delay_27_stateElements_6;
  reg        [254:0]  mulContext_delay_27_stateElements_7;
  reg        [254:0]  mulContext_delay_27_stateElements_8;
  reg        [254:0]  mulContext_delay_27_stateElements_9;
  reg        [254:0]  mulContext_delay_27_stateElements_10;
  reg                 mulContext_delay_28_isFull;
  reg        [2:0]    mulContext_delay_28_fullRound;
  reg        [5:0]    mulContext_delay_28_partialRound;
  reg        [3:0]    mulContext_delay_28_stateSize;
  reg        [7:0]    mulContext_delay_28_stateID;
  reg        [254:0]  mulContext_delay_28_stateElements_0;
  reg        [254:0]  mulContext_delay_28_stateElements_1;
  reg        [254:0]  mulContext_delay_28_stateElements_2;
  reg        [254:0]  mulContext_delay_28_stateElements_3;
  reg        [254:0]  mulContext_delay_28_stateElements_4;
  reg        [254:0]  mulContext_delay_28_stateElements_5;
  reg        [254:0]  mulContext_delay_28_stateElements_6;
  reg        [254:0]  mulContext_delay_28_stateElements_7;
  reg        [254:0]  mulContext_delay_28_stateElements_8;
  reg        [254:0]  mulContext_delay_28_stateElements_9;
  reg        [254:0]  mulContext_delay_28_stateElements_10;
  reg                 mulContext_delay_29_isFull;
  reg        [2:0]    mulContext_delay_29_fullRound;
  reg        [5:0]    mulContext_delay_29_partialRound;
  reg        [3:0]    mulContext_delay_29_stateSize;
  reg        [7:0]    mulContext_delay_29_stateID;
  reg        [254:0]  mulContext_delay_29_stateElements_0;
  reg        [254:0]  mulContext_delay_29_stateElements_1;
  reg        [254:0]  mulContext_delay_29_stateElements_2;
  reg        [254:0]  mulContext_delay_29_stateElements_3;
  reg        [254:0]  mulContext_delay_29_stateElements_4;
  reg        [254:0]  mulContext_delay_29_stateElements_5;
  reg        [254:0]  mulContext_delay_29_stateElements_6;
  reg        [254:0]  mulContext_delay_29_stateElements_7;
  reg        [254:0]  mulContext_delay_29_stateElements_8;
  reg        [254:0]  mulContext_delay_29_stateElements_9;
  reg        [254:0]  mulContext_delay_29_stateElements_10;
  reg                 mulContext_delay_30_isFull;
  reg        [2:0]    mulContext_delay_30_fullRound;
  reg        [5:0]    mulContext_delay_30_partialRound;
  reg        [3:0]    mulContext_delay_30_stateSize;
  reg        [7:0]    mulContext_delay_30_stateID;
  reg        [254:0]  mulContext_delay_30_stateElements_0;
  reg        [254:0]  mulContext_delay_30_stateElements_1;
  reg        [254:0]  mulContext_delay_30_stateElements_2;
  reg        [254:0]  mulContext_delay_30_stateElements_3;
  reg        [254:0]  mulContext_delay_30_stateElements_4;
  reg        [254:0]  mulContext_delay_30_stateElements_5;
  reg        [254:0]  mulContext_delay_30_stateElements_6;
  reg        [254:0]  mulContext_delay_30_stateElements_7;
  reg        [254:0]  mulContext_delay_30_stateElements_8;
  reg        [254:0]  mulContext_delay_30_stateElements_9;
  reg        [254:0]  mulContext_delay_30_stateElements_10;
  reg                 mulContext_delay_31_isFull;
  reg        [2:0]    mulContext_delay_31_fullRound;
  reg        [5:0]    mulContext_delay_31_partialRound;
  reg        [3:0]    mulContext_delay_31_stateSize;
  reg        [7:0]    mulContext_delay_31_stateID;
  reg        [254:0]  mulContext_delay_31_stateElements_0;
  reg        [254:0]  mulContext_delay_31_stateElements_1;
  reg        [254:0]  mulContext_delay_31_stateElements_2;
  reg        [254:0]  mulContext_delay_31_stateElements_3;
  reg        [254:0]  mulContext_delay_31_stateElements_4;
  reg        [254:0]  mulContext_delay_31_stateElements_5;
  reg        [254:0]  mulContext_delay_31_stateElements_6;
  reg        [254:0]  mulContext_delay_31_stateElements_7;
  reg        [254:0]  mulContext_delay_31_stateElements_8;
  reg        [254:0]  mulContext_delay_31_stateElements_9;
  reg        [254:0]  mulContext_delay_31_stateElements_10;
  reg                 mulContext_delay_32_isFull;
  reg        [2:0]    mulContext_delay_32_fullRound;
  reg        [5:0]    mulContext_delay_32_partialRound;
  reg        [3:0]    mulContext_delay_32_stateSize;
  reg        [7:0]    mulContext_delay_32_stateID;
  reg        [254:0]  mulContext_delay_32_stateElements_0;
  reg        [254:0]  mulContext_delay_32_stateElements_1;
  reg        [254:0]  mulContext_delay_32_stateElements_2;
  reg        [254:0]  mulContext_delay_32_stateElements_3;
  reg        [254:0]  mulContext_delay_32_stateElements_4;
  reg        [254:0]  mulContext_delay_32_stateElements_5;
  reg        [254:0]  mulContext_delay_32_stateElements_6;
  reg        [254:0]  mulContext_delay_32_stateElements_7;
  reg        [254:0]  mulContext_delay_32_stateElements_8;
  reg        [254:0]  mulContext_delay_32_stateElements_9;
  reg        [254:0]  mulContext_delay_32_stateElements_10;
  reg                 mulContext_delay_33_isFull;
  reg        [2:0]    mulContext_delay_33_fullRound;
  reg        [5:0]    mulContext_delay_33_partialRound;
  reg        [3:0]    mulContext_delay_33_stateSize;
  reg        [7:0]    mulContext_delay_33_stateID;
  reg        [254:0]  mulContext_delay_33_stateElements_0;
  reg        [254:0]  mulContext_delay_33_stateElements_1;
  reg        [254:0]  mulContext_delay_33_stateElements_2;
  reg        [254:0]  mulContext_delay_33_stateElements_3;
  reg        [254:0]  mulContext_delay_33_stateElements_4;
  reg        [254:0]  mulContext_delay_33_stateElements_5;
  reg        [254:0]  mulContext_delay_33_stateElements_6;
  reg        [254:0]  mulContext_delay_33_stateElements_7;
  reg        [254:0]  mulContext_delay_33_stateElements_8;
  reg        [254:0]  mulContext_delay_33_stateElements_9;
  reg        [254:0]  mulContext_delay_33_stateElements_10;
  reg                 mulContext_delay_34_isFull;
  reg        [2:0]    mulContext_delay_34_fullRound;
  reg        [5:0]    mulContext_delay_34_partialRound;
  reg        [3:0]    mulContext_delay_34_stateSize;
  reg        [7:0]    mulContext_delay_34_stateID;
  reg        [254:0]  mulContext_delay_34_stateElements_0;
  reg        [254:0]  mulContext_delay_34_stateElements_1;
  reg        [254:0]  mulContext_delay_34_stateElements_2;
  reg        [254:0]  mulContext_delay_34_stateElements_3;
  reg        [254:0]  mulContext_delay_34_stateElements_4;
  reg        [254:0]  mulContext_delay_34_stateElements_5;
  reg        [254:0]  mulContext_delay_34_stateElements_6;
  reg        [254:0]  mulContext_delay_34_stateElements_7;
  reg        [254:0]  mulContext_delay_34_stateElements_8;
  reg        [254:0]  mulContext_delay_34_stateElements_9;
  reg        [254:0]  mulContext_delay_34_stateElements_10;
  reg                 mulContext_delay_35_isFull;
  reg        [2:0]    mulContext_delay_35_fullRound;
  reg        [5:0]    mulContext_delay_35_partialRound;
  reg        [3:0]    mulContext_delay_35_stateSize;
  reg        [7:0]    mulContext_delay_35_stateID;
  reg        [254:0]  mulContext_delay_35_stateElements_0;
  reg        [254:0]  mulContext_delay_35_stateElements_1;
  reg        [254:0]  mulContext_delay_35_stateElements_2;
  reg        [254:0]  mulContext_delay_35_stateElements_3;
  reg        [254:0]  mulContext_delay_35_stateElements_4;
  reg        [254:0]  mulContext_delay_35_stateElements_5;
  reg        [254:0]  mulContext_delay_35_stateElements_6;
  reg        [254:0]  mulContext_delay_35_stateElements_7;
  reg        [254:0]  mulContext_delay_35_stateElements_8;
  reg        [254:0]  mulContext_delay_35_stateElements_9;
  reg        [254:0]  mulContext_delay_35_stateElements_10;
  reg                 mulContext_delay_36_isFull;
  reg        [2:0]    mulContext_delay_36_fullRound;
  reg        [5:0]    mulContext_delay_36_partialRound;
  reg        [3:0]    mulContext_delay_36_stateSize;
  reg        [7:0]    mulContext_delay_36_stateID;
  reg        [254:0]  mulContext_delay_36_stateElements_0;
  reg        [254:0]  mulContext_delay_36_stateElements_1;
  reg        [254:0]  mulContext_delay_36_stateElements_2;
  reg        [254:0]  mulContext_delay_36_stateElements_3;
  reg        [254:0]  mulContext_delay_36_stateElements_4;
  reg        [254:0]  mulContext_delay_36_stateElements_5;
  reg        [254:0]  mulContext_delay_36_stateElements_6;
  reg        [254:0]  mulContext_delay_36_stateElements_7;
  reg        [254:0]  mulContext_delay_36_stateElements_8;
  reg        [254:0]  mulContext_delay_36_stateElements_9;
  reg        [254:0]  mulContext_delay_36_stateElements_10;
  reg                 mulContext_delay_37_isFull;
  reg        [2:0]    mulContext_delay_37_fullRound;
  reg        [5:0]    mulContext_delay_37_partialRound;
  reg        [3:0]    mulContext_delay_37_stateSize;
  reg        [7:0]    mulContext_delay_37_stateID;
  reg        [254:0]  mulContext_delay_37_stateElements_0;
  reg        [254:0]  mulContext_delay_37_stateElements_1;
  reg        [254:0]  mulContext_delay_37_stateElements_2;
  reg        [254:0]  mulContext_delay_37_stateElements_3;
  reg        [254:0]  mulContext_delay_37_stateElements_4;
  reg        [254:0]  mulContext_delay_37_stateElements_5;
  reg        [254:0]  mulContext_delay_37_stateElements_6;
  reg        [254:0]  mulContext_delay_37_stateElements_7;
  reg        [254:0]  mulContext_delay_37_stateElements_8;
  reg        [254:0]  mulContext_delay_37_stateElements_9;
  reg        [254:0]  mulContext_delay_37_stateElements_10;
  reg                 mulContext_delay_38_isFull;
  reg        [2:0]    mulContext_delay_38_fullRound;
  reg        [5:0]    mulContext_delay_38_partialRound;
  reg        [3:0]    mulContext_delay_38_stateSize;
  reg        [7:0]    mulContext_delay_38_stateID;
  reg        [254:0]  mulContext_delay_38_stateElements_0;
  reg        [254:0]  mulContext_delay_38_stateElements_1;
  reg        [254:0]  mulContext_delay_38_stateElements_2;
  reg        [254:0]  mulContext_delay_38_stateElements_3;
  reg        [254:0]  mulContext_delay_38_stateElements_4;
  reg        [254:0]  mulContext_delay_38_stateElements_5;
  reg        [254:0]  mulContext_delay_38_stateElements_6;
  reg        [254:0]  mulContext_delay_38_stateElements_7;
  reg        [254:0]  mulContext_delay_38_stateElements_8;
  reg        [254:0]  mulContext_delay_38_stateElements_9;
  reg        [254:0]  mulContext_delay_38_stateElements_10;
  reg                 mulContext_delay_39_isFull;
  reg        [2:0]    mulContext_delay_39_fullRound;
  reg        [5:0]    mulContext_delay_39_partialRound;
  reg        [3:0]    mulContext_delay_39_stateSize;
  reg        [7:0]    mulContext_delay_39_stateID;
  reg        [254:0]  mulContext_delay_39_stateElements_0;
  reg        [254:0]  mulContext_delay_39_stateElements_1;
  reg        [254:0]  mulContext_delay_39_stateElements_2;
  reg        [254:0]  mulContext_delay_39_stateElements_3;
  reg        [254:0]  mulContext_delay_39_stateElements_4;
  reg        [254:0]  mulContext_delay_39_stateElements_5;
  reg        [254:0]  mulContext_delay_39_stateElements_6;
  reg        [254:0]  mulContext_delay_39_stateElements_7;
  reg        [254:0]  mulContext_delay_39_stateElements_8;
  reg        [254:0]  mulContext_delay_39_stateElements_9;
  reg        [254:0]  mulContext_delay_39_stateElements_10;
  reg                 mulContext_delay_40_isFull;
  reg        [2:0]    mulContext_delay_40_fullRound;
  reg        [5:0]    mulContext_delay_40_partialRound;
  reg        [3:0]    mulContext_delay_40_stateSize;
  reg        [7:0]    mulContext_delay_40_stateID;
  reg        [254:0]  mulContext_delay_40_stateElements_0;
  reg        [254:0]  mulContext_delay_40_stateElements_1;
  reg        [254:0]  mulContext_delay_40_stateElements_2;
  reg        [254:0]  mulContext_delay_40_stateElements_3;
  reg        [254:0]  mulContext_delay_40_stateElements_4;
  reg        [254:0]  mulContext_delay_40_stateElements_5;
  reg        [254:0]  mulContext_delay_40_stateElements_6;
  reg        [254:0]  mulContext_delay_40_stateElements_7;
  reg        [254:0]  mulContext_delay_40_stateElements_8;
  reg        [254:0]  mulContext_delay_40_stateElements_9;
  reg        [254:0]  mulContext_delay_40_stateElements_10;
  reg                 mulContext_delay_41_isFull;
  reg        [2:0]    mulContext_delay_41_fullRound;
  reg        [5:0]    mulContext_delay_41_partialRound;
  reg        [3:0]    mulContext_delay_41_stateSize;
  reg        [7:0]    mulContext_delay_41_stateID;
  reg        [254:0]  mulContext_delay_41_stateElements_0;
  reg        [254:0]  mulContext_delay_41_stateElements_1;
  reg        [254:0]  mulContext_delay_41_stateElements_2;
  reg        [254:0]  mulContext_delay_41_stateElements_3;
  reg        [254:0]  mulContext_delay_41_stateElements_4;
  reg        [254:0]  mulContext_delay_41_stateElements_5;
  reg        [254:0]  mulContext_delay_41_stateElements_6;
  reg        [254:0]  mulContext_delay_41_stateElements_7;
  reg        [254:0]  mulContext_delay_41_stateElements_8;
  reg        [254:0]  mulContext_delay_41_stateElements_9;
  reg        [254:0]  mulContext_delay_41_stateElements_10;
  reg                 mulContext_delay_42_isFull;
  reg        [2:0]    mulContext_delay_42_fullRound;
  reg        [5:0]    mulContext_delay_42_partialRound;
  reg        [3:0]    mulContext_delay_42_stateSize;
  reg        [7:0]    mulContext_delay_42_stateID;
  reg        [254:0]  mulContext_delay_42_stateElements_0;
  reg        [254:0]  mulContext_delay_42_stateElements_1;
  reg        [254:0]  mulContext_delay_42_stateElements_2;
  reg        [254:0]  mulContext_delay_42_stateElements_3;
  reg        [254:0]  mulContext_delay_42_stateElements_4;
  reg        [254:0]  mulContext_delay_42_stateElements_5;
  reg        [254:0]  mulContext_delay_42_stateElements_6;
  reg        [254:0]  mulContext_delay_42_stateElements_7;
  reg        [254:0]  mulContext_delay_42_stateElements_8;
  reg        [254:0]  mulContext_delay_42_stateElements_9;
  reg        [254:0]  mulContext_delay_42_stateElements_10;
  reg                 mulContext_delay_43_isFull;
  reg        [2:0]    mulContext_delay_43_fullRound;
  reg        [5:0]    mulContext_delay_43_partialRound;
  reg        [3:0]    mulContext_delay_43_stateSize;
  reg        [7:0]    mulContext_delay_43_stateID;
  reg        [254:0]  mulContext_delay_43_stateElements_0;
  reg        [254:0]  mulContext_delay_43_stateElements_1;
  reg        [254:0]  mulContext_delay_43_stateElements_2;
  reg        [254:0]  mulContext_delay_43_stateElements_3;
  reg        [254:0]  mulContext_delay_43_stateElements_4;
  reg        [254:0]  mulContext_delay_43_stateElements_5;
  reg        [254:0]  mulContext_delay_43_stateElements_6;
  reg        [254:0]  mulContext_delay_43_stateElements_7;
  reg        [254:0]  mulContext_delay_43_stateElements_8;
  reg        [254:0]  mulContext_delay_43_stateElements_9;
  reg        [254:0]  mulContext_delay_43_stateElements_10;
  reg                 mulContext_delay_44_isFull;
  reg        [2:0]    mulContext_delay_44_fullRound;
  reg        [5:0]    mulContext_delay_44_partialRound;
  reg        [3:0]    mulContext_delay_44_stateSize;
  reg        [7:0]    mulContext_delay_44_stateID;
  reg        [254:0]  mulContext_delay_44_stateElements_0;
  reg        [254:0]  mulContext_delay_44_stateElements_1;
  reg        [254:0]  mulContext_delay_44_stateElements_2;
  reg        [254:0]  mulContext_delay_44_stateElements_3;
  reg        [254:0]  mulContext_delay_44_stateElements_4;
  reg        [254:0]  mulContext_delay_44_stateElements_5;
  reg        [254:0]  mulContext_delay_44_stateElements_6;
  reg        [254:0]  mulContext_delay_44_stateElements_7;
  reg        [254:0]  mulContext_delay_44_stateElements_8;
  reg        [254:0]  mulContext_delay_44_stateElements_9;
  reg        [254:0]  mulContext_delay_44_stateElements_10;
  reg                 mulContext_delay_45_isFull;
  reg        [2:0]    mulContext_delay_45_fullRound;
  reg        [5:0]    mulContext_delay_45_partialRound;
  reg        [3:0]    mulContext_delay_45_stateSize;
  reg        [7:0]    mulContext_delay_45_stateID;
  reg        [254:0]  mulContext_delay_45_stateElements_0;
  reg        [254:0]  mulContext_delay_45_stateElements_1;
  reg        [254:0]  mulContext_delay_45_stateElements_2;
  reg        [254:0]  mulContext_delay_45_stateElements_3;
  reg        [254:0]  mulContext_delay_45_stateElements_4;
  reg        [254:0]  mulContext_delay_45_stateElements_5;
  reg        [254:0]  mulContext_delay_45_stateElements_6;
  reg        [254:0]  mulContext_delay_45_stateElements_7;
  reg        [254:0]  mulContext_delay_45_stateElements_8;
  reg        [254:0]  mulContext_delay_45_stateElements_9;
  reg        [254:0]  mulContext_delay_45_stateElements_10;
  reg                 mulContext_delay_46_isFull;
  reg        [2:0]    mulContext_delay_46_fullRound;
  reg        [5:0]    mulContext_delay_46_partialRound;
  reg        [3:0]    mulContext_delay_46_stateSize;
  reg        [7:0]    mulContext_delay_46_stateID;
  reg        [254:0]  mulContext_delay_46_stateElements_0;
  reg        [254:0]  mulContext_delay_46_stateElements_1;
  reg        [254:0]  mulContext_delay_46_stateElements_2;
  reg        [254:0]  mulContext_delay_46_stateElements_3;
  reg        [254:0]  mulContext_delay_46_stateElements_4;
  reg        [254:0]  mulContext_delay_46_stateElements_5;
  reg        [254:0]  mulContext_delay_46_stateElements_6;
  reg        [254:0]  mulContext_delay_46_stateElements_7;
  reg        [254:0]  mulContext_delay_46_stateElements_8;
  reg        [254:0]  mulContext_delay_46_stateElements_9;
  reg        [254:0]  mulContext_delay_46_stateElements_10;
  reg                 mulContext_delay_47_isFull;
  reg        [2:0]    mulContext_delay_47_fullRound;
  reg        [5:0]    mulContext_delay_47_partialRound;
  reg        [3:0]    mulContext_delay_47_stateSize;
  reg        [7:0]    mulContext_delay_47_stateID;
  reg        [254:0]  mulContext_delay_47_stateElements_0;
  reg        [254:0]  mulContext_delay_47_stateElements_1;
  reg        [254:0]  mulContext_delay_47_stateElements_2;
  reg        [254:0]  mulContext_delay_47_stateElements_3;
  reg        [254:0]  mulContext_delay_47_stateElements_4;
  reg        [254:0]  mulContext_delay_47_stateElements_5;
  reg        [254:0]  mulContext_delay_47_stateElements_6;
  reg        [254:0]  mulContext_delay_47_stateElements_7;
  reg        [254:0]  mulContext_delay_47_stateElements_8;
  reg        [254:0]  mulContext_delay_47_stateElements_9;
  reg        [254:0]  mulContext_delay_47_stateElements_10;
  reg                 mulContext_delay_48_isFull;
  reg        [2:0]    mulContext_delay_48_fullRound;
  reg        [5:0]    mulContext_delay_48_partialRound;
  reg        [3:0]    mulContext_delay_48_stateSize;
  reg        [7:0]    mulContext_delay_48_stateID;
  reg        [254:0]  mulContext_delay_48_stateElements_0;
  reg        [254:0]  mulContext_delay_48_stateElements_1;
  reg        [254:0]  mulContext_delay_48_stateElements_2;
  reg        [254:0]  mulContext_delay_48_stateElements_3;
  reg        [254:0]  mulContext_delay_48_stateElements_4;
  reg        [254:0]  mulContext_delay_48_stateElements_5;
  reg        [254:0]  mulContext_delay_48_stateElements_6;
  reg        [254:0]  mulContext_delay_48_stateElements_7;
  reg        [254:0]  mulContext_delay_48_stateElements_8;
  reg        [254:0]  mulContext_delay_48_stateElements_9;
  reg        [254:0]  mulContext_delay_48_stateElements_10;
  reg                 mulContext_delay_49_isFull;
  reg        [2:0]    mulContext_delay_49_fullRound;
  reg        [5:0]    mulContext_delay_49_partialRound;
  reg        [3:0]    mulContext_delay_49_stateSize;
  reg        [7:0]    mulContext_delay_49_stateID;
  reg        [254:0]  mulContext_delay_49_stateElements_0;
  reg        [254:0]  mulContext_delay_49_stateElements_1;
  reg        [254:0]  mulContext_delay_49_stateElements_2;
  reg        [254:0]  mulContext_delay_49_stateElements_3;
  reg        [254:0]  mulContext_delay_49_stateElements_4;
  reg        [254:0]  mulContext_delay_49_stateElements_5;
  reg        [254:0]  mulContext_delay_49_stateElements_6;
  reg        [254:0]  mulContext_delay_49_stateElements_7;
  reg        [254:0]  mulContext_delay_49_stateElements_8;
  reg        [254:0]  mulContext_delay_49_stateElements_9;
  reg        [254:0]  mulContext_delay_49_stateElements_10;
  reg                 mulContextDelayed_isFull;
  reg        [2:0]    mulContextDelayed_fullRound;
  reg        [5:0]    mulContextDelayed_partialRound;
  reg        [3:0]    mulContextDelayed_stateSize;
  reg        [7:0]    mulContextDelayed_stateID;
  reg        [254:0]  mulContextDelayed_stateElements_0;
  reg        [254:0]  mulContextDelayed_stateElements_1;
  reg        [254:0]  mulContextDelayed_stateElements_2;
  reg        [254:0]  mulContextDelayed_stateElements_3;
  reg        [254:0]  mulContextDelayed_stateElements_4;
  reg        [254:0]  mulContextDelayed_stateElements_5;
  reg        [254:0]  mulContextDelayed_stateElements_6;
  reg        [254:0]  mulContextDelayed_stateElements_7;
  reg        [254:0]  mulContextDelayed_stateElements_8;
  reg        [254:0]  mulContextDelayed_stateElements_9;
  reg        [254:0]  mulContextDelayed_stateElements_10;
  reg                 _zz_validDelayed;
  reg                 _zz_validDelayed_1;
  reg                 _zz_validDelayed_2;
  reg                 _zz_validDelayed_3;
  reg                 _zz_validDelayed_4;
  reg                 _zz_validDelayed_5;
  reg                 _zz_validDelayed_6;
  reg                 _zz_validDelayed_7;
  reg                 _zz_validDelayed_8;
  reg                 _zz_validDelayed_9;
  reg                 _zz_validDelayed_10;
  reg                 _zz_validDelayed_11;
  reg                 _zz_validDelayed_12;
  reg                 _zz_validDelayed_13;
  reg                 _zz_validDelayed_14;
  reg                 validDelayed;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_1;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_2;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_3;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_4;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_5;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_6;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_7;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_8;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_9;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_10;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_11;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_12;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_13;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_14;
  reg        [254:0]  montgomeryMultFlow_15_io_output_payload_res_delay_15;
  reg        [254:0]  mulOutput0Delayed;
  wire                addContext_isFull;
  wire       [2:0]    addContext_fullRound;
  wire       [5:0]    addContext_partialRound;
  wire       [3:0]    addContext_stateSize;
  wire       [7:0]    addContext_stateID;
  reg                 addContext_delay_1_isFull;
  reg        [2:0]    addContext_delay_1_fullRound;
  reg        [5:0]    addContext_delay_1_partialRound;
  reg        [3:0]    addContext_delay_1_stateSize;
  reg        [7:0]    addContext_delay_1_stateID;
  reg                 addContext_delay_2_isFull;
  reg        [2:0]    addContext_delay_2_fullRound;
  reg        [5:0]    addContext_delay_2_partialRound;
  reg        [3:0]    addContext_delay_2_stateSize;
  reg        [7:0]    addContext_delay_2_stateID;
  reg                 addContext_delay_3_isFull;
  reg        [2:0]    addContext_delay_3_fullRound;
  reg        [5:0]    addContext_delay_3_partialRound;
  reg        [3:0]    addContext_delay_3_stateSize;
  reg        [7:0]    addContext_delay_3_stateID;
  reg                 addContext_delay_4_isFull;
  reg        [2:0]    addContext_delay_4_fullRound;
  reg        [5:0]    addContext_delay_4_partialRound;
  reg        [3:0]    addContext_delay_4_stateSize;
  reg        [7:0]    addContext_delay_4_stateID;
  reg                 addContext_delay_5_isFull;
  reg        [2:0]    addContext_delay_5_fullRound;
  reg        [5:0]    addContext_delay_5_partialRound;
  reg        [3:0]    addContext_delay_5_stateSize;
  reg        [7:0]    addContext_delay_5_stateID;
  reg                 addContext_delay_6_isFull;
  reg        [2:0]    addContext_delay_6_fullRound;
  reg        [5:0]    addContext_delay_6_partialRound;
  reg        [3:0]    addContext_delay_6_stateSize;
  reg        [7:0]    addContext_delay_6_stateID;
  reg                 addContext_delay_7_isFull;
  reg        [2:0]    addContext_delay_7_fullRound;
  reg        [5:0]    addContext_delay_7_partialRound;
  reg        [3:0]    addContext_delay_7_stateSize;
  reg        [7:0]    addContext_delay_7_stateID;
  reg                 addContext_delay_8_isFull;
  reg        [2:0]    addContext_delay_8_fullRound;
  reg        [5:0]    addContext_delay_8_partialRound;
  reg        [3:0]    addContext_delay_8_stateSize;
  reg        [7:0]    addContext_delay_8_stateID;
  reg                 addContext_delay_9_isFull;
  reg        [2:0]    addContext_delay_9_fullRound;
  reg        [5:0]    addContext_delay_9_partialRound;
  reg        [3:0]    addContext_delay_9_stateSize;
  reg        [7:0]    addContext_delay_9_stateID;
  reg                 addContext_delay_10_isFull;
  reg        [2:0]    addContext_delay_10_fullRound;
  reg        [5:0]    addContext_delay_10_partialRound;
  reg        [3:0]    addContext_delay_10_stateSize;
  reg        [7:0]    addContext_delay_10_stateID;
  reg                 addContext_delay_11_isFull;
  reg        [2:0]    addContext_delay_11_fullRound;
  reg        [5:0]    addContext_delay_11_partialRound;
  reg        [3:0]    addContext_delay_11_stateSize;
  reg        [7:0]    addContext_delay_11_stateID;
  reg                 addContext_delay_12_isFull;
  reg        [2:0]    addContext_delay_12_fullRound;
  reg        [5:0]    addContext_delay_12_partialRound;
  reg        [3:0]    addContext_delay_12_stateSize;
  reg        [7:0]    addContext_delay_12_stateID;
  reg                 addContext_delay_13_isFull;
  reg        [2:0]    addContext_delay_13_fullRound;
  reg        [5:0]    addContext_delay_13_partialRound;
  reg        [3:0]    addContext_delay_13_stateSize;
  reg        [7:0]    addContext_delay_13_stateID;
  reg                 addContext_delay_14_isFull;
  reg        [2:0]    addContext_delay_14_fullRound;
  reg        [5:0]    addContext_delay_14_partialRound;
  reg        [3:0]    addContext_delay_14_stateSize;
  reg        [7:0]    addContext_delay_14_stateID;
  reg                 addContext_delay_15_isFull;
  reg        [2:0]    addContext_delay_15_fullRound;
  reg        [5:0]    addContext_delay_15_partialRound;
  reg        [3:0]    addContext_delay_15_stateSize;
  reg        [7:0]    addContext_delay_15_stateID;
  reg                 addContextDelayed_isFull;
  reg        [2:0]    addContextDelayed_fullRound;
  reg        [5:0]    addContextDelayed_partialRound;
  reg        [3:0]    addContextDelayed_stateSize;
  reg        [7:0]    addContextDelayed_stateID;
  wire       [3059:0] _zz_io_output_payload_stateElements_0;

  assign _zz__zz_validDelayed = montgomeryMultFlow_16_io_output_valid;
  assign _zz__zz_validDelayed_1 = montgomeryMultFlow_15_io_output_valid;
  assign _zz__zz_io_output_payload_stateElements_0 = modAdderPiped_23_io_res;
  assign _zz__zz_io_output_payload_stateElements_0_1 = modAdderPiped_22_io_res;
  MDSConstantMem constants (
    .io_addr_isFull          (io_input_payload_isFull             ), //i
    .io_addr_fullRound       (io_input_payload_fullRound[2:0]     ), //i
    .io_addr_partialRound    (io_input_payload_partialRound[5:0]  ), //i
    .io_addr_stateIndex      (io_input_payload_stateIndex[3:0]    ), //i
    .io_addr_stateSize       (io_input_payload_stateSize[3:0]     ), //i
    .io_data_0               (constants_io_data_0[254:0]          ), //o
    .io_data_1               (constants_io_data_1[254:0]          ), //o
    .io_data_2               (constants_io_data_2[254:0]          ), //o
    .io_data_3               (constants_io_data_3[254:0]          ), //o
    .io_data_4               (constants_io_data_4[254:0]          ), //o
    .io_data_5               (constants_io_data_5[254:0]          ), //o
    .io_data_6               (constants_io_data_6[254:0]          ), //o
    .io_data_7               (constants_io_data_7[254:0]          ), //o
    .io_data_8               (constants_io_data_8[254:0]          ), //o
    .io_data_9               (constants_io_data_9[254:0]          ), //o
    .io_data_10              (constants_io_data_10[254:0]         ), //o
    .io_data_11              (constants_io_data_11[254:0]         ), //o
    .clk                     (clk                                 ), //i
    .resetn                  (resetn                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_15 (
    .io_input_valid           (mulInputsTemp_0_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_0_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_0_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_15_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_15_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_16 (
    .io_input_valid           (mulInputsTemp_1_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_1_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_1_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_16_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_16_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_17 (
    .io_input_valid           (mulInputsTemp_2_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_2_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_2_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_17_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_17_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_18 (
    .io_input_valid           (mulInputsTemp_3_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_3_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_3_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_18_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_18_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_19 (
    .io_input_valid           (mulInputsTemp_4_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_4_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_4_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_19_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_19_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_20 (
    .io_input_valid           (mulInputsTemp_5_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_5_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_5_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_20_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_20_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_21 (
    .io_input_valid           (mulInputsTemp_6_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_6_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_6_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_21_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_21_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_22 (
    .io_input_valid           (mulInputsTemp_7_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_7_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_7_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_22_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_22_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_23 (
    .io_input_valid           (mulInputsTemp_8_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_8_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_8_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_23_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_23_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_24 (
    .io_input_valid           (mulInputsTemp_9_valid                               ), //i
    .io_input_payload_op1     (mulInputsTemp_9_payload_op1[254:0]                  ), //i
    .io_input_payload_op2     (mulInputsTemp_9_payload_op2[254:0]                  ), //i
    .io_output_valid          (montgomeryMultFlow_24_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_24_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_25 (
    .io_input_valid           (mulInputsTemp_10_valid                              ), //i
    .io_input_payload_op1     (mulInputsTemp_10_payload_op1[254:0]                 ), //i
    .io_input_payload_op2     (mulInputsTemp_10_payload_op2[254:0]                 ), //i
    .io_output_valid          (montgomeryMultFlow_25_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_25_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  MontgomeryMultFlow montgomeryMultFlow_26 (
    .io_input_valid           (mulInputsTemp_11_valid                              ), //i
    .io_input_payload_op1     (mulInputsTemp_11_payload_op1[254:0]                 ), //i
    .io_input_payload_op2     (mulInputsTemp_11_payload_op2[254:0]                 ), //i
    .io_output_valid          (montgomeryMultFlow_26_io_output_valid               ), //o
    .io_output_payload_res    (montgomeryMultFlow_26_io_output_payload_res[254:0]  ), //o
    .clk                      (clk                                                 ), //i
    .resetn                   (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_22 (
    .io_op1    (montgomeryMultFlow_16_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_0[254:0]            ), //i
    .io_res    (modAdderPiped_22_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_23 (
    .io_op1    (montgomeryMultFlow_17_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_1[254:0]            ), //i
    .io_res    (modAdderPiped_23_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_24 (
    .io_op1    (montgomeryMultFlow_18_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_2[254:0]            ), //i
    .io_res    (modAdderPiped_24_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_25 (
    .io_op1    (montgomeryMultFlow_19_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_3[254:0]            ), //i
    .io_res    (modAdderPiped_25_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_26 (
    .io_op1    (montgomeryMultFlow_20_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_4[254:0]            ), //i
    .io_res    (modAdderPiped_26_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_27 (
    .io_op1    (montgomeryMultFlow_21_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_5[254:0]            ), //i
    .io_res    (modAdderPiped_27_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_28 (
    .io_op1    (montgomeryMultFlow_22_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_6[254:0]            ), //i
    .io_res    (modAdderPiped_28_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_29 (
    .io_op1    (montgomeryMultFlow_23_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_7[254:0]            ), //i
    .io_res    (modAdderPiped_29_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_30 (
    .io_op1    (montgomeryMultFlow_24_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_8[254:0]            ), //i
    .io_res    (modAdderPiped_30_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_31 (
    .io_op1    (montgomeryMultFlow_25_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_9[254:0]            ), //i
    .io_res    (modAdderPiped_31_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  ModAdderPiped modAdderPiped_32 (
    .io_op1    (montgomeryMultFlow_26_io_output_payload_res[254:0]  ), //i
    .io_op2    (mulContextDelayed_stateElements_10[254:0]           ), //i
    .io_res    (modAdderPiped_32_io_res[254:0]                      ), //o
    .clk       (clk                                                 ), //i
    .resetn    (resetn                                              )  //i
  );
  assign mulInputs_0_valid = inputDelayed_valid;
  assign mulInputs_0_payload_op1 = inputDelayed_payload_stateElement;
  assign mulInputs_0_payload_op2 = constants_io_data_0;
  assign mulInputs_1_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_1_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(!when_MDSMatrixMultiplier_l74) begin
        if(!when_MDSMatrixMultiplier_l76) begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_1_payload_op1 = inputDelayed_payload_stateElements_0;
          end
        end
      end
    end
  end

  assign mulInputs_1_payload_op2 = constants_io_data_1;
  assign mulInputs_2_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_2_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(!when_MDSMatrixMultiplier_l74) begin
        if(!when_MDSMatrixMultiplier_l76) begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_2_payload_op1 = inputDelayed_payload_stateElements_1;
          end
        end
      end
    end
  end

  assign mulInputs_2_payload_op2 = constants_io_data_2;
  assign mulInputs_3_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_3_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(when_MDSMatrixMultiplier_l74) begin
        mulInputs_3_payload_op1 = inputDelayed_payload_stateElements_0;
      end else begin
        if(!when_MDSMatrixMultiplier_l76) begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_3_payload_op1 = inputDelayed_payload_stateElements_2;
          end
        end
      end
    end
  end

  assign mulInputs_3_payload_op2 = constants_io_data_3;
  assign mulInputs_4_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_4_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(when_MDSMatrixMultiplier_l74) begin
        mulInputs_4_payload_op1 = inputDelayed_payload_stateElements_1;
      end else begin
        if(!when_MDSMatrixMultiplier_l76) begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_4_payload_op1 = inputDelayed_payload_stateElements_3;
          end
        end
      end
    end
  end

  assign mulInputs_4_payload_op2 = constants_io_data_4;
  assign mulInputs_5_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_5_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(!when_MDSMatrixMultiplier_l74) begin
        if(when_MDSMatrixMultiplier_l76) begin
          mulInputs_5_payload_op1 = inputDelayed_payload_stateElements_0;
        end else begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_5_payload_op1 = inputDelayed_payload_stateElements_4;
          end
        end
      end
    end
  end

  assign mulInputs_5_payload_op2 = constants_io_data_5;
  assign mulInputs_6_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_6_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(!when_MDSMatrixMultiplier_l74) begin
        if(when_MDSMatrixMultiplier_l76) begin
          mulInputs_6_payload_op1 = inputDelayed_payload_stateElements_1;
        end else begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_6_payload_op1 = inputDelayed_payload_stateElements_5;
          end
        end
      end
    end
  end

  assign mulInputs_6_payload_op2 = constants_io_data_6;
  assign mulInputs_7_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_7_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(!when_MDSMatrixMultiplier_l74) begin
        if(when_MDSMatrixMultiplier_l76) begin
          mulInputs_7_payload_op1 = inputDelayed_payload_stateElements_2;
        end else begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_7_payload_op1 = inputDelayed_payload_stateElements_6;
          end
        end
      end
    end
  end

  assign mulInputs_7_payload_op2 = constants_io_data_7;
  assign mulInputs_8_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_8_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(!when_MDSMatrixMultiplier_l74) begin
        if(when_MDSMatrixMultiplier_l76) begin
          mulInputs_8_payload_op1 = inputDelayed_payload_stateElements_3;
        end else begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_8_payload_op1 = inputDelayed_payload_stateElements_7;
          end
        end
      end
    end
  end

  assign mulInputs_8_payload_op2 = constants_io_data_8;
  assign mulInputs_9_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_9_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(!when_MDSMatrixMultiplier_l74) begin
        if(!when_MDSMatrixMultiplier_l76) begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_9_payload_op1 = inputDelayed_payload_stateElements_8;
          end
        end
      end
    end
  end

  assign mulInputs_9_payload_op2 = constants_io_data_9;
  assign mulInputs_10_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_10_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(!when_MDSMatrixMultiplier_l74) begin
        if(!when_MDSMatrixMultiplier_l76) begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_10_payload_op1 = inputDelayed_payload_stateElements_9;
          end
        end
      end
    end
  end

  assign mulInputs_10_payload_op2 = constants_io_data_10;
  assign mulInputs_11_valid = inputDelayed_valid;
  always @(*) begin
    mulInputs_11_payload_op1 = inputDelayed_payload_stateElement;
    if(when_MDSMatrixMultiplier_l73) begin
      if(!when_MDSMatrixMultiplier_l74) begin
        if(!when_MDSMatrixMultiplier_l76) begin
          if(when_MDSMatrixMultiplier_l78) begin
            mulInputs_11_payload_op1 = inputDelayed_payload_stateElements_10;
          end
        end
      end
    end
  end

  assign mulInputs_11_payload_op2 = constants_io_data_11;
  assign when_MDSMatrixMultiplier_l73 = (! inputDelayed_payload_isFull);
  assign when_MDSMatrixMultiplier_l74 = (inputDelayed_payload_stateSize == 4'b0011);
  assign when_MDSMatrixMultiplier_l76 = (inputDelayed_payload_stateSize == 4'b0101);
  assign when_MDSMatrixMultiplier_l78 = (inputDelayed_payload_stateIndex == 4'b0001);
  assign mulContext_isFull = inputDelayed_payload_isFull;
  assign mulContext_fullRound = inputDelayed_payload_fullRound;
  assign mulContext_partialRound = inputDelayed_payload_partialRound;
  assign mulContext_stateSize = inputDelayed_payload_stateSize;
  assign mulContext_stateID = inputDelayed_payload_stateID;
  always @(*) begin
    mulContext_stateElements_0 = inputDelayed_payload_stateElements_0;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_0 = _zz_mulContext_stateElements_0[254 : 0];
    end
  end

  always @(*) begin
    mulContext_stateElements_1 = inputDelayed_payload_stateElements_1;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_1 = _zz_mulContext_stateElements_0[509 : 255];
    end
  end

  always @(*) begin
    mulContext_stateElements_2 = inputDelayed_payload_stateElements_2;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_2 = _zz_mulContext_stateElements_0[764 : 510];
    end
  end

  always @(*) begin
    mulContext_stateElements_3 = inputDelayed_payload_stateElements_3;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_3 = _zz_mulContext_stateElements_0[1019 : 765];
    end
  end

  always @(*) begin
    mulContext_stateElements_4 = inputDelayed_payload_stateElements_4;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_4 = _zz_mulContext_stateElements_0[1274 : 1020];
    end
  end

  always @(*) begin
    mulContext_stateElements_5 = inputDelayed_payload_stateElements_5;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_5 = _zz_mulContext_stateElements_0[1529 : 1275];
    end
  end

  always @(*) begin
    mulContext_stateElements_6 = inputDelayed_payload_stateElements_6;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_6 = _zz_mulContext_stateElements_0[1784 : 1530];
    end
  end

  always @(*) begin
    mulContext_stateElements_7 = inputDelayed_payload_stateElements_7;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_7 = _zz_mulContext_stateElements_0[2039 : 1785];
    end
  end

  always @(*) begin
    mulContext_stateElements_8 = inputDelayed_payload_stateElements_8;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_8 = _zz_mulContext_stateElements_0[2294 : 2040];
    end
  end

  always @(*) begin
    mulContext_stateElements_9 = inputDelayed_payload_stateElements_9;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_9 = _zz_mulContext_stateElements_0[2549 : 2295];
    end
  end

  always @(*) begin
    mulContext_stateElements_10 = inputDelayed_payload_stateElements_10;
    if(when_MDSMatrixMultiplier_l94) begin
      mulContext_stateElements_10 = _zz_mulContext_stateElements_0[2804 : 2550];
    end
  end

  assign when_MDSMatrixMultiplier_l94 = (((! inputDelayed_payload_isFull) && (4'b0101 < inputDelayed_payload_stateSize)) && (inputDelayed_payload_stateIndex == 4'b0001));
  assign _zz_mulContext_stateElements_0 = 2805'h0;
  assign addContext_isFull = mulContextDelayed_isFull;
  assign addContext_fullRound = mulContextDelayed_fullRound;
  assign addContext_partialRound = mulContextDelayed_partialRound;
  assign addContext_stateSize = mulContextDelayed_stateSize;
  assign addContext_stateID = mulContextDelayed_stateID;
  assign io_output_valid = validDelayed;
  assign io_output_payload_isFull = addContextDelayed_isFull;
  assign io_output_payload_fullRound = addContextDelayed_fullRound;
  assign io_output_payload_partialRound = addContextDelayed_partialRound;
  assign io_output_payload_stateSize = addContextDelayed_stateSize;
  assign io_output_payload_stateID = addContextDelayed_stateID;
  assign _zz_io_output_payload_stateElements_0 = {{modAdderPiped_32_io_res,{modAdderPiped_31_io_res,{modAdderPiped_30_io_res,{modAdderPiped_29_io_res,{modAdderPiped_28_io_res,{modAdderPiped_27_io_res,{modAdderPiped_26_io_res,{modAdderPiped_25_io_res,{modAdderPiped_24_io_res,{_zz__zz_io_output_payload_stateElements_0,_zz__zz_io_output_payload_stateElements_0_1}}}}}}}}}},mulOutput0Delayed};
  assign io_output_payload_stateElements_0 = _zz_io_output_payload_stateElements_0[254 : 0];
  assign io_output_payload_stateElements_1 = _zz_io_output_payload_stateElements_0[509 : 255];
  assign io_output_payload_stateElements_2 = _zz_io_output_payload_stateElements_0[764 : 510];
  assign io_output_payload_stateElements_3 = _zz_io_output_payload_stateElements_0[1019 : 765];
  assign io_output_payload_stateElements_4 = _zz_io_output_payload_stateElements_0[1274 : 1020];
  assign io_output_payload_stateElements_5 = _zz_io_output_payload_stateElements_0[1529 : 1275];
  assign io_output_payload_stateElements_6 = _zz_io_output_payload_stateElements_0[1784 : 1530];
  assign io_output_payload_stateElements_7 = _zz_io_output_payload_stateElements_0[2039 : 1785];
  assign io_output_payload_stateElements_8 = _zz_io_output_payload_stateElements_0[2294 : 2040];
  assign io_output_payload_stateElements_9 = _zz_io_output_payload_stateElements_0[2549 : 2295];
  assign io_output_payload_stateElements_10 = _zz_io_output_payload_stateElements_0[2804 : 2550];
  assign io_output_payload_stateElements_11 = _zz_io_output_payload_stateElements_0[3059 : 2805];
  always @(posedge clk) begin
    if(!resetn) begin
      io_input_regNext_valid <= 1'b0;
      io_input_regNext_regNext_valid <= 1'b0;
      io_input_regNext_regNext_regNext_valid <= 1'b0;
      io_input_regNext_regNext_regNext_regNext_valid <= 1'b0;
      inputDelayed_valid <= 1'b0;
      mulInputsTemp_0_valid <= 1'b0;
      mulInputsTemp_1_valid <= 1'b0;
      mulInputsTemp_2_valid <= 1'b0;
      mulInputsTemp_3_valid <= 1'b0;
      mulInputsTemp_4_valid <= 1'b0;
      mulInputsTemp_5_valid <= 1'b0;
      mulInputsTemp_6_valid <= 1'b0;
      mulInputsTemp_7_valid <= 1'b0;
      mulInputsTemp_8_valid <= 1'b0;
      mulInputsTemp_9_valid <= 1'b0;
      mulInputsTemp_10_valid <= 1'b0;
      mulInputsTemp_11_valid <= 1'b0;
      _zz_validDelayed <= 1'b0;
      _zz_validDelayed_1 <= 1'b0;
      _zz_validDelayed_2 <= 1'b0;
      _zz_validDelayed_3 <= 1'b0;
      _zz_validDelayed_4 <= 1'b0;
      _zz_validDelayed_5 <= 1'b0;
      _zz_validDelayed_6 <= 1'b0;
      _zz_validDelayed_7 <= 1'b0;
      _zz_validDelayed_8 <= 1'b0;
      _zz_validDelayed_9 <= 1'b0;
      _zz_validDelayed_10 <= 1'b0;
      _zz_validDelayed_11 <= 1'b0;
      _zz_validDelayed_12 <= 1'b0;
      _zz_validDelayed_13 <= 1'b0;
      _zz_validDelayed_14 <= 1'b0;
      validDelayed <= 1'b0;
    end else begin
      io_input_regNext_valid <= io_input_valid;
      io_input_regNext_regNext_valid <= io_input_regNext_valid;
      io_input_regNext_regNext_regNext_valid <= io_input_regNext_regNext_valid;
      io_input_regNext_regNext_regNext_regNext_valid <= io_input_regNext_regNext_regNext_valid;
      inputDelayed_valid <= io_input_regNext_regNext_regNext_regNext_valid;
      mulInputsTemp_0_valid <= mulInputs_0_valid;
      mulInputsTemp_1_valid <= mulInputs_1_valid;
      mulInputsTemp_2_valid <= mulInputs_2_valid;
      mulInputsTemp_3_valid <= mulInputs_3_valid;
      mulInputsTemp_4_valid <= mulInputs_4_valid;
      mulInputsTemp_5_valid <= mulInputs_5_valid;
      mulInputsTemp_6_valid <= mulInputs_6_valid;
      mulInputsTemp_7_valid <= mulInputs_7_valid;
      mulInputsTemp_8_valid <= mulInputs_8_valid;
      mulInputsTemp_9_valid <= mulInputs_9_valid;
      mulInputsTemp_10_valid <= mulInputs_10_valid;
      mulInputsTemp_11_valid <= mulInputs_11_valid;
      _zz_validDelayed <= (&{montgomeryMultFlow_26_io_output_valid,{montgomeryMultFlow_25_io_output_valid,{montgomeryMultFlow_24_io_output_valid,{montgomeryMultFlow_23_io_output_valid,{montgomeryMultFlow_22_io_output_valid,{montgomeryMultFlow_21_io_output_valid,{montgomeryMultFlow_20_io_output_valid,{montgomeryMultFlow_19_io_output_valid,{montgomeryMultFlow_18_io_output_valid,{montgomeryMultFlow_17_io_output_valid,{_zz__zz_validDelayed,_zz__zz_validDelayed_1}}}}}}}}}}});
      _zz_validDelayed_1 <= _zz_validDelayed;
      _zz_validDelayed_2 <= _zz_validDelayed_1;
      _zz_validDelayed_3 <= _zz_validDelayed_2;
      _zz_validDelayed_4 <= _zz_validDelayed_3;
      _zz_validDelayed_5 <= _zz_validDelayed_4;
      _zz_validDelayed_6 <= _zz_validDelayed_5;
      _zz_validDelayed_7 <= _zz_validDelayed_6;
      _zz_validDelayed_8 <= _zz_validDelayed_7;
      _zz_validDelayed_9 <= _zz_validDelayed_8;
      _zz_validDelayed_10 <= _zz_validDelayed_9;
      _zz_validDelayed_11 <= _zz_validDelayed_10;
      _zz_validDelayed_12 <= _zz_validDelayed_11;
      _zz_validDelayed_13 <= _zz_validDelayed_12;
      _zz_validDelayed_14 <= _zz_validDelayed_13;
      validDelayed <= _zz_validDelayed_14;
    end
  end

  always @(posedge clk) begin
    io_input_regNext_payload_isFull <= io_input_payload_isFull;
    io_input_regNext_payload_fullRound <= io_input_payload_fullRound;
    io_input_regNext_payload_partialRound <= io_input_payload_partialRound;
    io_input_regNext_payload_stateIndex <= io_input_payload_stateIndex;
    io_input_regNext_payload_stateSize <= io_input_payload_stateSize;
    io_input_regNext_payload_stateID <= io_input_payload_stateID;
    io_input_regNext_payload_stateElements_0 <= io_input_payload_stateElements_0;
    io_input_regNext_payload_stateElements_1 <= io_input_payload_stateElements_1;
    io_input_regNext_payload_stateElements_2 <= io_input_payload_stateElements_2;
    io_input_regNext_payload_stateElements_3 <= io_input_payload_stateElements_3;
    io_input_regNext_payload_stateElements_4 <= io_input_payload_stateElements_4;
    io_input_regNext_payload_stateElements_5 <= io_input_payload_stateElements_5;
    io_input_regNext_payload_stateElements_6 <= io_input_payload_stateElements_6;
    io_input_regNext_payload_stateElements_7 <= io_input_payload_stateElements_7;
    io_input_regNext_payload_stateElements_8 <= io_input_payload_stateElements_8;
    io_input_regNext_payload_stateElements_9 <= io_input_payload_stateElements_9;
    io_input_regNext_payload_stateElements_10 <= io_input_payload_stateElements_10;
    io_input_regNext_payload_stateElement <= io_input_payload_stateElement;
    io_input_regNext_regNext_payload_isFull <= io_input_regNext_payload_isFull;
    io_input_regNext_regNext_payload_fullRound <= io_input_regNext_payload_fullRound;
    io_input_regNext_regNext_payload_partialRound <= io_input_regNext_payload_partialRound;
    io_input_regNext_regNext_payload_stateIndex <= io_input_regNext_payload_stateIndex;
    io_input_regNext_regNext_payload_stateSize <= io_input_regNext_payload_stateSize;
    io_input_regNext_regNext_payload_stateID <= io_input_regNext_payload_stateID;
    io_input_regNext_regNext_payload_stateElements_0 <= io_input_regNext_payload_stateElements_0;
    io_input_regNext_regNext_payload_stateElements_1 <= io_input_regNext_payload_stateElements_1;
    io_input_regNext_regNext_payload_stateElements_2 <= io_input_regNext_payload_stateElements_2;
    io_input_regNext_regNext_payload_stateElements_3 <= io_input_regNext_payload_stateElements_3;
    io_input_regNext_regNext_payload_stateElements_4 <= io_input_regNext_payload_stateElements_4;
    io_input_regNext_regNext_payload_stateElements_5 <= io_input_regNext_payload_stateElements_5;
    io_input_regNext_regNext_payload_stateElements_6 <= io_input_regNext_payload_stateElements_6;
    io_input_regNext_regNext_payload_stateElements_7 <= io_input_regNext_payload_stateElements_7;
    io_input_regNext_regNext_payload_stateElements_8 <= io_input_regNext_payload_stateElements_8;
    io_input_regNext_regNext_payload_stateElements_9 <= io_input_regNext_payload_stateElements_9;
    io_input_regNext_regNext_payload_stateElements_10 <= io_input_regNext_payload_stateElements_10;
    io_input_regNext_regNext_payload_stateElement <= io_input_regNext_payload_stateElement;
    io_input_regNext_regNext_regNext_payload_isFull <= io_input_regNext_regNext_payload_isFull;
    io_input_regNext_regNext_regNext_payload_fullRound <= io_input_regNext_regNext_payload_fullRound;
    io_input_regNext_regNext_regNext_payload_partialRound <= io_input_regNext_regNext_payload_partialRound;
    io_input_regNext_regNext_regNext_payload_stateIndex <= io_input_regNext_regNext_payload_stateIndex;
    io_input_regNext_regNext_regNext_payload_stateSize <= io_input_regNext_regNext_payload_stateSize;
    io_input_regNext_regNext_regNext_payload_stateID <= io_input_regNext_regNext_payload_stateID;
    io_input_regNext_regNext_regNext_payload_stateElements_0 <= io_input_regNext_regNext_payload_stateElements_0;
    io_input_regNext_regNext_regNext_payload_stateElements_1 <= io_input_regNext_regNext_payload_stateElements_1;
    io_input_regNext_regNext_regNext_payload_stateElements_2 <= io_input_regNext_regNext_payload_stateElements_2;
    io_input_regNext_regNext_regNext_payload_stateElements_3 <= io_input_regNext_regNext_payload_stateElements_3;
    io_input_regNext_regNext_regNext_payload_stateElements_4 <= io_input_regNext_regNext_payload_stateElements_4;
    io_input_regNext_regNext_regNext_payload_stateElements_5 <= io_input_regNext_regNext_payload_stateElements_5;
    io_input_regNext_regNext_regNext_payload_stateElements_6 <= io_input_regNext_regNext_payload_stateElements_6;
    io_input_regNext_regNext_regNext_payload_stateElements_7 <= io_input_regNext_regNext_payload_stateElements_7;
    io_input_regNext_regNext_regNext_payload_stateElements_8 <= io_input_regNext_regNext_payload_stateElements_8;
    io_input_regNext_regNext_regNext_payload_stateElements_9 <= io_input_regNext_regNext_payload_stateElements_9;
    io_input_regNext_regNext_regNext_payload_stateElements_10 <= io_input_regNext_regNext_payload_stateElements_10;
    io_input_regNext_regNext_regNext_payload_stateElement <= io_input_regNext_regNext_payload_stateElement;
    io_input_regNext_regNext_regNext_regNext_payload_isFull <= io_input_regNext_regNext_regNext_payload_isFull;
    io_input_regNext_regNext_regNext_regNext_payload_fullRound <= io_input_regNext_regNext_regNext_payload_fullRound;
    io_input_regNext_regNext_regNext_regNext_payload_partialRound <= io_input_regNext_regNext_regNext_payload_partialRound;
    io_input_regNext_regNext_regNext_regNext_payload_stateIndex <= io_input_regNext_regNext_regNext_payload_stateIndex;
    io_input_regNext_regNext_regNext_regNext_payload_stateSize <= io_input_regNext_regNext_regNext_payload_stateSize;
    io_input_regNext_regNext_regNext_regNext_payload_stateID <= io_input_regNext_regNext_regNext_payload_stateID;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_0 <= io_input_regNext_regNext_regNext_payload_stateElements_0;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_1 <= io_input_regNext_regNext_regNext_payload_stateElements_1;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_2 <= io_input_regNext_regNext_regNext_payload_stateElements_2;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_3 <= io_input_regNext_regNext_regNext_payload_stateElements_3;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_4 <= io_input_regNext_regNext_regNext_payload_stateElements_4;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_5 <= io_input_regNext_regNext_regNext_payload_stateElements_5;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_6 <= io_input_regNext_regNext_regNext_payload_stateElements_6;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_7 <= io_input_regNext_regNext_regNext_payload_stateElements_7;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_8 <= io_input_regNext_regNext_regNext_payload_stateElements_8;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_9 <= io_input_regNext_regNext_regNext_payload_stateElements_9;
    io_input_regNext_regNext_regNext_regNext_payload_stateElements_10 <= io_input_regNext_regNext_regNext_payload_stateElements_10;
    io_input_regNext_regNext_regNext_regNext_payload_stateElement <= io_input_regNext_regNext_regNext_payload_stateElement;
    inputDelayed_payload_isFull <= io_input_regNext_regNext_regNext_regNext_payload_isFull;
    inputDelayed_payload_fullRound <= io_input_regNext_regNext_regNext_regNext_payload_fullRound;
    inputDelayed_payload_partialRound <= io_input_regNext_regNext_regNext_regNext_payload_partialRound;
    inputDelayed_payload_stateIndex <= io_input_regNext_regNext_regNext_regNext_payload_stateIndex;
    inputDelayed_payload_stateSize <= io_input_regNext_regNext_regNext_regNext_payload_stateSize;
    inputDelayed_payload_stateID <= io_input_regNext_regNext_regNext_regNext_payload_stateID;
    inputDelayed_payload_stateElements_0 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_0;
    inputDelayed_payload_stateElements_1 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_1;
    inputDelayed_payload_stateElements_2 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_2;
    inputDelayed_payload_stateElements_3 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_3;
    inputDelayed_payload_stateElements_4 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_4;
    inputDelayed_payload_stateElements_5 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_5;
    inputDelayed_payload_stateElements_6 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_6;
    inputDelayed_payload_stateElements_7 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_7;
    inputDelayed_payload_stateElements_8 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_8;
    inputDelayed_payload_stateElements_9 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_9;
    inputDelayed_payload_stateElements_10 <= io_input_regNext_regNext_regNext_regNext_payload_stateElements_10;
    inputDelayed_payload_stateElement <= io_input_regNext_regNext_regNext_regNext_payload_stateElement;
    mulInputsTemp_0_payload_op1 <= mulInputs_0_payload_op1;
    mulInputsTemp_0_payload_op2 <= mulInputs_0_payload_op2;
    mulInputsTemp_1_payload_op1 <= mulInputs_1_payload_op1;
    mulInputsTemp_1_payload_op2 <= mulInputs_1_payload_op2;
    mulInputsTemp_2_payload_op1 <= mulInputs_2_payload_op1;
    mulInputsTemp_2_payload_op2 <= mulInputs_2_payload_op2;
    mulInputsTemp_3_payload_op1 <= mulInputs_3_payload_op1;
    mulInputsTemp_3_payload_op2 <= mulInputs_3_payload_op2;
    mulInputsTemp_4_payload_op1 <= mulInputs_4_payload_op1;
    mulInputsTemp_4_payload_op2 <= mulInputs_4_payload_op2;
    mulInputsTemp_5_payload_op1 <= mulInputs_5_payload_op1;
    mulInputsTemp_5_payload_op2 <= mulInputs_5_payload_op2;
    mulInputsTemp_6_payload_op1 <= mulInputs_6_payload_op1;
    mulInputsTemp_6_payload_op2 <= mulInputs_6_payload_op2;
    mulInputsTemp_7_payload_op1 <= mulInputs_7_payload_op1;
    mulInputsTemp_7_payload_op2 <= mulInputs_7_payload_op2;
    mulInputsTemp_8_payload_op1 <= mulInputs_8_payload_op1;
    mulInputsTemp_8_payload_op2 <= mulInputs_8_payload_op2;
    mulInputsTemp_9_payload_op1 <= mulInputs_9_payload_op1;
    mulInputsTemp_9_payload_op2 <= mulInputs_9_payload_op2;
    mulInputsTemp_10_payload_op1 <= mulInputs_10_payload_op1;
    mulInputsTemp_10_payload_op2 <= mulInputs_10_payload_op2;
    mulInputsTemp_11_payload_op1 <= mulInputs_11_payload_op1;
    mulInputsTemp_11_payload_op2 <= mulInputs_11_payload_op2;
    mulContext_delay_1_isFull <= mulContext_isFull;
    mulContext_delay_1_fullRound <= mulContext_fullRound;
    mulContext_delay_1_partialRound <= mulContext_partialRound;
    mulContext_delay_1_stateSize <= mulContext_stateSize;
    mulContext_delay_1_stateID <= mulContext_stateID;
    mulContext_delay_1_stateElements_0 <= mulContext_stateElements_0;
    mulContext_delay_1_stateElements_1 <= mulContext_stateElements_1;
    mulContext_delay_1_stateElements_2 <= mulContext_stateElements_2;
    mulContext_delay_1_stateElements_3 <= mulContext_stateElements_3;
    mulContext_delay_1_stateElements_4 <= mulContext_stateElements_4;
    mulContext_delay_1_stateElements_5 <= mulContext_stateElements_5;
    mulContext_delay_1_stateElements_6 <= mulContext_stateElements_6;
    mulContext_delay_1_stateElements_7 <= mulContext_stateElements_7;
    mulContext_delay_1_stateElements_8 <= mulContext_stateElements_8;
    mulContext_delay_1_stateElements_9 <= mulContext_stateElements_9;
    mulContext_delay_1_stateElements_10 <= mulContext_stateElements_10;
    mulContext_delay_2_isFull <= mulContext_delay_1_isFull;
    mulContext_delay_2_fullRound <= mulContext_delay_1_fullRound;
    mulContext_delay_2_partialRound <= mulContext_delay_1_partialRound;
    mulContext_delay_2_stateSize <= mulContext_delay_1_stateSize;
    mulContext_delay_2_stateID <= mulContext_delay_1_stateID;
    mulContext_delay_2_stateElements_0 <= mulContext_delay_1_stateElements_0;
    mulContext_delay_2_stateElements_1 <= mulContext_delay_1_stateElements_1;
    mulContext_delay_2_stateElements_2 <= mulContext_delay_1_stateElements_2;
    mulContext_delay_2_stateElements_3 <= mulContext_delay_1_stateElements_3;
    mulContext_delay_2_stateElements_4 <= mulContext_delay_1_stateElements_4;
    mulContext_delay_2_stateElements_5 <= mulContext_delay_1_stateElements_5;
    mulContext_delay_2_stateElements_6 <= mulContext_delay_1_stateElements_6;
    mulContext_delay_2_stateElements_7 <= mulContext_delay_1_stateElements_7;
    mulContext_delay_2_stateElements_8 <= mulContext_delay_1_stateElements_8;
    mulContext_delay_2_stateElements_9 <= mulContext_delay_1_stateElements_9;
    mulContext_delay_2_stateElements_10 <= mulContext_delay_1_stateElements_10;
    mulContext_delay_3_isFull <= mulContext_delay_2_isFull;
    mulContext_delay_3_fullRound <= mulContext_delay_2_fullRound;
    mulContext_delay_3_partialRound <= mulContext_delay_2_partialRound;
    mulContext_delay_3_stateSize <= mulContext_delay_2_stateSize;
    mulContext_delay_3_stateID <= mulContext_delay_2_stateID;
    mulContext_delay_3_stateElements_0 <= mulContext_delay_2_stateElements_0;
    mulContext_delay_3_stateElements_1 <= mulContext_delay_2_stateElements_1;
    mulContext_delay_3_stateElements_2 <= mulContext_delay_2_stateElements_2;
    mulContext_delay_3_stateElements_3 <= mulContext_delay_2_stateElements_3;
    mulContext_delay_3_stateElements_4 <= mulContext_delay_2_stateElements_4;
    mulContext_delay_3_stateElements_5 <= mulContext_delay_2_stateElements_5;
    mulContext_delay_3_stateElements_6 <= mulContext_delay_2_stateElements_6;
    mulContext_delay_3_stateElements_7 <= mulContext_delay_2_stateElements_7;
    mulContext_delay_3_stateElements_8 <= mulContext_delay_2_stateElements_8;
    mulContext_delay_3_stateElements_9 <= mulContext_delay_2_stateElements_9;
    mulContext_delay_3_stateElements_10 <= mulContext_delay_2_stateElements_10;
    mulContext_delay_4_isFull <= mulContext_delay_3_isFull;
    mulContext_delay_4_fullRound <= mulContext_delay_3_fullRound;
    mulContext_delay_4_partialRound <= mulContext_delay_3_partialRound;
    mulContext_delay_4_stateSize <= mulContext_delay_3_stateSize;
    mulContext_delay_4_stateID <= mulContext_delay_3_stateID;
    mulContext_delay_4_stateElements_0 <= mulContext_delay_3_stateElements_0;
    mulContext_delay_4_stateElements_1 <= mulContext_delay_3_stateElements_1;
    mulContext_delay_4_stateElements_2 <= mulContext_delay_3_stateElements_2;
    mulContext_delay_4_stateElements_3 <= mulContext_delay_3_stateElements_3;
    mulContext_delay_4_stateElements_4 <= mulContext_delay_3_stateElements_4;
    mulContext_delay_4_stateElements_5 <= mulContext_delay_3_stateElements_5;
    mulContext_delay_4_stateElements_6 <= mulContext_delay_3_stateElements_6;
    mulContext_delay_4_stateElements_7 <= mulContext_delay_3_stateElements_7;
    mulContext_delay_4_stateElements_8 <= mulContext_delay_3_stateElements_8;
    mulContext_delay_4_stateElements_9 <= mulContext_delay_3_stateElements_9;
    mulContext_delay_4_stateElements_10 <= mulContext_delay_3_stateElements_10;
    mulContext_delay_5_isFull <= mulContext_delay_4_isFull;
    mulContext_delay_5_fullRound <= mulContext_delay_4_fullRound;
    mulContext_delay_5_partialRound <= mulContext_delay_4_partialRound;
    mulContext_delay_5_stateSize <= mulContext_delay_4_stateSize;
    mulContext_delay_5_stateID <= mulContext_delay_4_stateID;
    mulContext_delay_5_stateElements_0 <= mulContext_delay_4_stateElements_0;
    mulContext_delay_5_stateElements_1 <= mulContext_delay_4_stateElements_1;
    mulContext_delay_5_stateElements_2 <= mulContext_delay_4_stateElements_2;
    mulContext_delay_5_stateElements_3 <= mulContext_delay_4_stateElements_3;
    mulContext_delay_5_stateElements_4 <= mulContext_delay_4_stateElements_4;
    mulContext_delay_5_stateElements_5 <= mulContext_delay_4_stateElements_5;
    mulContext_delay_5_stateElements_6 <= mulContext_delay_4_stateElements_6;
    mulContext_delay_5_stateElements_7 <= mulContext_delay_4_stateElements_7;
    mulContext_delay_5_stateElements_8 <= mulContext_delay_4_stateElements_8;
    mulContext_delay_5_stateElements_9 <= mulContext_delay_4_stateElements_9;
    mulContext_delay_5_stateElements_10 <= mulContext_delay_4_stateElements_10;
    mulContext_delay_6_isFull <= mulContext_delay_5_isFull;
    mulContext_delay_6_fullRound <= mulContext_delay_5_fullRound;
    mulContext_delay_6_partialRound <= mulContext_delay_5_partialRound;
    mulContext_delay_6_stateSize <= mulContext_delay_5_stateSize;
    mulContext_delay_6_stateID <= mulContext_delay_5_stateID;
    mulContext_delay_6_stateElements_0 <= mulContext_delay_5_stateElements_0;
    mulContext_delay_6_stateElements_1 <= mulContext_delay_5_stateElements_1;
    mulContext_delay_6_stateElements_2 <= mulContext_delay_5_stateElements_2;
    mulContext_delay_6_stateElements_3 <= mulContext_delay_5_stateElements_3;
    mulContext_delay_6_stateElements_4 <= mulContext_delay_5_stateElements_4;
    mulContext_delay_6_stateElements_5 <= mulContext_delay_5_stateElements_5;
    mulContext_delay_6_stateElements_6 <= mulContext_delay_5_stateElements_6;
    mulContext_delay_6_stateElements_7 <= mulContext_delay_5_stateElements_7;
    mulContext_delay_6_stateElements_8 <= mulContext_delay_5_stateElements_8;
    mulContext_delay_6_stateElements_9 <= mulContext_delay_5_stateElements_9;
    mulContext_delay_6_stateElements_10 <= mulContext_delay_5_stateElements_10;
    mulContext_delay_7_isFull <= mulContext_delay_6_isFull;
    mulContext_delay_7_fullRound <= mulContext_delay_6_fullRound;
    mulContext_delay_7_partialRound <= mulContext_delay_6_partialRound;
    mulContext_delay_7_stateSize <= mulContext_delay_6_stateSize;
    mulContext_delay_7_stateID <= mulContext_delay_6_stateID;
    mulContext_delay_7_stateElements_0 <= mulContext_delay_6_stateElements_0;
    mulContext_delay_7_stateElements_1 <= mulContext_delay_6_stateElements_1;
    mulContext_delay_7_stateElements_2 <= mulContext_delay_6_stateElements_2;
    mulContext_delay_7_stateElements_3 <= mulContext_delay_6_stateElements_3;
    mulContext_delay_7_stateElements_4 <= mulContext_delay_6_stateElements_4;
    mulContext_delay_7_stateElements_5 <= mulContext_delay_6_stateElements_5;
    mulContext_delay_7_stateElements_6 <= mulContext_delay_6_stateElements_6;
    mulContext_delay_7_stateElements_7 <= mulContext_delay_6_stateElements_7;
    mulContext_delay_7_stateElements_8 <= mulContext_delay_6_stateElements_8;
    mulContext_delay_7_stateElements_9 <= mulContext_delay_6_stateElements_9;
    mulContext_delay_7_stateElements_10 <= mulContext_delay_6_stateElements_10;
    mulContext_delay_8_isFull <= mulContext_delay_7_isFull;
    mulContext_delay_8_fullRound <= mulContext_delay_7_fullRound;
    mulContext_delay_8_partialRound <= mulContext_delay_7_partialRound;
    mulContext_delay_8_stateSize <= mulContext_delay_7_stateSize;
    mulContext_delay_8_stateID <= mulContext_delay_7_stateID;
    mulContext_delay_8_stateElements_0 <= mulContext_delay_7_stateElements_0;
    mulContext_delay_8_stateElements_1 <= mulContext_delay_7_stateElements_1;
    mulContext_delay_8_stateElements_2 <= mulContext_delay_7_stateElements_2;
    mulContext_delay_8_stateElements_3 <= mulContext_delay_7_stateElements_3;
    mulContext_delay_8_stateElements_4 <= mulContext_delay_7_stateElements_4;
    mulContext_delay_8_stateElements_5 <= mulContext_delay_7_stateElements_5;
    mulContext_delay_8_stateElements_6 <= mulContext_delay_7_stateElements_6;
    mulContext_delay_8_stateElements_7 <= mulContext_delay_7_stateElements_7;
    mulContext_delay_8_stateElements_8 <= mulContext_delay_7_stateElements_8;
    mulContext_delay_8_stateElements_9 <= mulContext_delay_7_stateElements_9;
    mulContext_delay_8_stateElements_10 <= mulContext_delay_7_stateElements_10;
    mulContext_delay_9_isFull <= mulContext_delay_8_isFull;
    mulContext_delay_9_fullRound <= mulContext_delay_8_fullRound;
    mulContext_delay_9_partialRound <= mulContext_delay_8_partialRound;
    mulContext_delay_9_stateSize <= mulContext_delay_8_stateSize;
    mulContext_delay_9_stateID <= mulContext_delay_8_stateID;
    mulContext_delay_9_stateElements_0 <= mulContext_delay_8_stateElements_0;
    mulContext_delay_9_stateElements_1 <= mulContext_delay_8_stateElements_1;
    mulContext_delay_9_stateElements_2 <= mulContext_delay_8_stateElements_2;
    mulContext_delay_9_stateElements_3 <= mulContext_delay_8_stateElements_3;
    mulContext_delay_9_stateElements_4 <= mulContext_delay_8_stateElements_4;
    mulContext_delay_9_stateElements_5 <= mulContext_delay_8_stateElements_5;
    mulContext_delay_9_stateElements_6 <= mulContext_delay_8_stateElements_6;
    mulContext_delay_9_stateElements_7 <= mulContext_delay_8_stateElements_7;
    mulContext_delay_9_stateElements_8 <= mulContext_delay_8_stateElements_8;
    mulContext_delay_9_stateElements_9 <= mulContext_delay_8_stateElements_9;
    mulContext_delay_9_stateElements_10 <= mulContext_delay_8_stateElements_10;
    mulContext_delay_10_isFull <= mulContext_delay_9_isFull;
    mulContext_delay_10_fullRound <= mulContext_delay_9_fullRound;
    mulContext_delay_10_partialRound <= mulContext_delay_9_partialRound;
    mulContext_delay_10_stateSize <= mulContext_delay_9_stateSize;
    mulContext_delay_10_stateID <= mulContext_delay_9_stateID;
    mulContext_delay_10_stateElements_0 <= mulContext_delay_9_stateElements_0;
    mulContext_delay_10_stateElements_1 <= mulContext_delay_9_stateElements_1;
    mulContext_delay_10_stateElements_2 <= mulContext_delay_9_stateElements_2;
    mulContext_delay_10_stateElements_3 <= mulContext_delay_9_stateElements_3;
    mulContext_delay_10_stateElements_4 <= mulContext_delay_9_stateElements_4;
    mulContext_delay_10_stateElements_5 <= mulContext_delay_9_stateElements_5;
    mulContext_delay_10_stateElements_6 <= mulContext_delay_9_stateElements_6;
    mulContext_delay_10_stateElements_7 <= mulContext_delay_9_stateElements_7;
    mulContext_delay_10_stateElements_8 <= mulContext_delay_9_stateElements_8;
    mulContext_delay_10_stateElements_9 <= mulContext_delay_9_stateElements_9;
    mulContext_delay_10_stateElements_10 <= mulContext_delay_9_stateElements_10;
    mulContext_delay_11_isFull <= mulContext_delay_10_isFull;
    mulContext_delay_11_fullRound <= mulContext_delay_10_fullRound;
    mulContext_delay_11_partialRound <= mulContext_delay_10_partialRound;
    mulContext_delay_11_stateSize <= mulContext_delay_10_stateSize;
    mulContext_delay_11_stateID <= mulContext_delay_10_stateID;
    mulContext_delay_11_stateElements_0 <= mulContext_delay_10_stateElements_0;
    mulContext_delay_11_stateElements_1 <= mulContext_delay_10_stateElements_1;
    mulContext_delay_11_stateElements_2 <= mulContext_delay_10_stateElements_2;
    mulContext_delay_11_stateElements_3 <= mulContext_delay_10_stateElements_3;
    mulContext_delay_11_stateElements_4 <= mulContext_delay_10_stateElements_4;
    mulContext_delay_11_stateElements_5 <= mulContext_delay_10_stateElements_5;
    mulContext_delay_11_stateElements_6 <= mulContext_delay_10_stateElements_6;
    mulContext_delay_11_stateElements_7 <= mulContext_delay_10_stateElements_7;
    mulContext_delay_11_stateElements_8 <= mulContext_delay_10_stateElements_8;
    mulContext_delay_11_stateElements_9 <= mulContext_delay_10_stateElements_9;
    mulContext_delay_11_stateElements_10 <= mulContext_delay_10_stateElements_10;
    mulContext_delay_12_isFull <= mulContext_delay_11_isFull;
    mulContext_delay_12_fullRound <= mulContext_delay_11_fullRound;
    mulContext_delay_12_partialRound <= mulContext_delay_11_partialRound;
    mulContext_delay_12_stateSize <= mulContext_delay_11_stateSize;
    mulContext_delay_12_stateID <= mulContext_delay_11_stateID;
    mulContext_delay_12_stateElements_0 <= mulContext_delay_11_stateElements_0;
    mulContext_delay_12_stateElements_1 <= mulContext_delay_11_stateElements_1;
    mulContext_delay_12_stateElements_2 <= mulContext_delay_11_stateElements_2;
    mulContext_delay_12_stateElements_3 <= mulContext_delay_11_stateElements_3;
    mulContext_delay_12_stateElements_4 <= mulContext_delay_11_stateElements_4;
    mulContext_delay_12_stateElements_5 <= mulContext_delay_11_stateElements_5;
    mulContext_delay_12_stateElements_6 <= mulContext_delay_11_stateElements_6;
    mulContext_delay_12_stateElements_7 <= mulContext_delay_11_stateElements_7;
    mulContext_delay_12_stateElements_8 <= mulContext_delay_11_stateElements_8;
    mulContext_delay_12_stateElements_9 <= mulContext_delay_11_stateElements_9;
    mulContext_delay_12_stateElements_10 <= mulContext_delay_11_stateElements_10;
    mulContext_delay_13_isFull <= mulContext_delay_12_isFull;
    mulContext_delay_13_fullRound <= mulContext_delay_12_fullRound;
    mulContext_delay_13_partialRound <= mulContext_delay_12_partialRound;
    mulContext_delay_13_stateSize <= mulContext_delay_12_stateSize;
    mulContext_delay_13_stateID <= mulContext_delay_12_stateID;
    mulContext_delay_13_stateElements_0 <= mulContext_delay_12_stateElements_0;
    mulContext_delay_13_stateElements_1 <= mulContext_delay_12_stateElements_1;
    mulContext_delay_13_stateElements_2 <= mulContext_delay_12_stateElements_2;
    mulContext_delay_13_stateElements_3 <= mulContext_delay_12_stateElements_3;
    mulContext_delay_13_stateElements_4 <= mulContext_delay_12_stateElements_4;
    mulContext_delay_13_stateElements_5 <= mulContext_delay_12_stateElements_5;
    mulContext_delay_13_stateElements_6 <= mulContext_delay_12_stateElements_6;
    mulContext_delay_13_stateElements_7 <= mulContext_delay_12_stateElements_7;
    mulContext_delay_13_stateElements_8 <= mulContext_delay_12_stateElements_8;
    mulContext_delay_13_stateElements_9 <= mulContext_delay_12_stateElements_9;
    mulContext_delay_13_stateElements_10 <= mulContext_delay_12_stateElements_10;
    mulContext_delay_14_isFull <= mulContext_delay_13_isFull;
    mulContext_delay_14_fullRound <= mulContext_delay_13_fullRound;
    mulContext_delay_14_partialRound <= mulContext_delay_13_partialRound;
    mulContext_delay_14_stateSize <= mulContext_delay_13_stateSize;
    mulContext_delay_14_stateID <= mulContext_delay_13_stateID;
    mulContext_delay_14_stateElements_0 <= mulContext_delay_13_stateElements_0;
    mulContext_delay_14_stateElements_1 <= mulContext_delay_13_stateElements_1;
    mulContext_delay_14_stateElements_2 <= mulContext_delay_13_stateElements_2;
    mulContext_delay_14_stateElements_3 <= mulContext_delay_13_stateElements_3;
    mulContext_delay_14_stateElements_4 <= mulContext_delay_13_stateElements_4;
    mulContext_delay_14_stateElements_5 <= mulContext_delay_13_stateElements_5;
    mulContext_delay_14_stateElements_6 <= mulContext_delay_13_stateElements_6;
    mulContext_delay_14_stateElements_7 <= mulContext_delay_13_stateElements_7;
    mulContext_delay_14_stateElements_8 <= mulContext_delay_13_stateElements_8;
    mulContext_delay_14_stateElements_9 <= mulContext_delay_13_stateElements_9;
    mulContext_delay_14_stateElements_10 <= mulContext_delay_13_stateElements_10;
    mulContext_delay_15_isFull <= mulContext_delay_14_isFull;
    mulContext_delay_15_fullRound <= mulContext_delay_14_fullRound;
    mulContext_delay_15_partialRound <= mulContext_delay_14_partialRound;
    mulContext_delay_15_stateSize <= mulContext_delay_14_stateSize;
    mulContext_delay_15_stateID <= mulContext_delay_14_stateID;
    mulContext_delay_15_stateElements_0 <= mulContext_delay_14_stateElements_0;
    mulContext_delay_15_stateElements_1 <= mulContext_delay_14_stateElements_1;
    mulContext_delay_15_stateElements_2 <= mulContext_delay_14_stateElements_2;
    mulContext_delay_15_stateElements_3 <= mulContext_delay_14_stateElements_3;
    mulContext_delay_15_stateElements_4 <= mulContext_delay_14_stateElements_4;
    mulContext_delay_15_stateElements_5 <= mulContext_delay_14_stateElements_5;
    mulContext_delay_15_stateElements_6 <= mulContext_delay_14_stateElements_6;
    mulContext_delay_15_stateElements_7 <= mulContext_delay_14_stateElements_7;
    mulContext_delay_15_stateElements_8 <= mulContext_delay_14_stateElements_8;
    mulContext_delay_15_stateElements_9 <= mulContext_delay_14_stateElements_9;
    mulContext_delay_15_stateElements_10 <= mulContext_delay_14_stateElements_10;
    mulContext_delay_16_isFull <= mulContext_delay_15_isFull;
    mulContext_delay_16_fullRound <= mulContext_delay_15_fullRound;
    mulContext_delay_16_partialRound <= mulContext_delay_15_partialRound;
    mulContext_delay_16_stateSize <= mulContext_delay_15_stateSize;
    mulContext_delay_16_stateID <= mulContext_delay_15_stateID;
    mulContext_delay_16_stateElements_0 <= mulContext_delay_15_stateElements_0;
    mulContext_delay_16_stateElements_1 <= mulContext_delay_15_stateElements_1;
    mulContext_delay_16_stateElements_2 <= mulContext_delay_15_stateElements_2;
    mulContext_delay_16_stateElements_3 <= mulContext_delay_15_stateElements_3;
    mulContext_delay_16_stateElements_4 <= mulContext_delay_15_stateElements_4;
    mulContext_delay_16_stateElements_5 <= mulContext_delay_15_stateElements_5;
    mulContext_delay_16_stateElements_6 <= mulContext_delay_15_stateElements_6;
    mulContext_delay_16_stateElements_7 <= mulContext_delay_15_stateElements_7;
    mulContext_delay_16_stateElements_8 <= mulContext_delay_15_stateElements_8;
    mulContext_delay_16_stateElements_9 <= mulContext_delay_15_stateElements_9;
    mulContext_delay_16_stateElements_10 <= mulContext_delay_15_stateElements_10;
    mulContext_delay_17_isFull <= mulContext_delay_16_isFull;
    mulContext_delay_17_fullRound <= mulContext_delay_16_fullRound;
    mulContext_delay_17_partialRound <= mulContext_delay_16_partialRound;
    mulContext_delay_17_stateSize <= mulContext_delay_16_stateSize;
    mulContext_delay_17_stateID <= mulContext_delay_16_stateID;
    mulContext_delay_17_stateElements_0 <= mulContext_delay_16_stateElements_0;
    mulContext_delay_17_stateElements_1 <= mulContext_delay_16_stateElements_1;
    mulContext_delay_17_stateElements_2 <= mulContext_delay_16_stateElements_2;
    mulContext_delay_17_stateElements_3 <= mulContext_delay_16_stateElements_3;
    mulContext_delay_17_stateElements_4 <= mulContext_delay_16_stateElements_4;
    mulContext_delay_17_stateElements_5 <= mulContext_delay_16_stateElements_5;
    mulContext_delay_17_stateElements_6 <= mulContext_delay_16_stateElements_6;
    mulContext_delay_17_stateElements_7 <= mulContext_delay_16_stateElements_7;
    mulContext_delay_17_stateElements_8 <= mulContext_delay_16_stateElements_8;
    mulContext_delay_17_stateElements_9 <= mulContext_delay_16_stateElements_9;
    mulContext_delay_17_stateElements_10 <= mulContext_delay_16_stateElements_10;
    mulContext_delay_18_isFull <= mulContext_delay_17_isFull;
    mulContext_delay_18_fullRound <= mulContext_delay_17_fullRound;
    mulContext_delay_18_partialRound <= mulContext_delay_17_partialRound;
    mulContext_delay_18_stateSize <= mulContext_delay_17_stateSize;
    mulContext_delay_18_stateID <= mulContext_delay_17_stateID;
    mulContext_delay_18_stateElements_0 <= mulContext_delay_17_stateElements_0;
    mulContext_delay_18_stateElements_1 <= mulContext_delay_17_stateElements_1;
    mulContext_delay_18_stateElements_2 <= mulContext_delay_17_stateElements_2;
    mulContext_delay_18_stateElements_3 <= mulContext_delay_17_stateElements_3;
    mulContext_delay_18_stateElements_4 <= mulContext_delay_17_stateElements_4;
    mulContext_delay_18_stateElements_5 <= mulContext_delay_17_stateElements_5;
    mulContext_delay_18_stateElements_6 <= mulContext_delay_17_stateElements_6;
    mulContext_delay_18_stateElements_7 <= mulContext_delay_17_stateElements_7;
    mulContext_delay_18_stateElements_8 <= mulContext_delay_17_stateElements_8;
    mulContext_delay_18_stateElements_9 <= mulContext_delay_17_stateElements_9;
    mulContext_delay_18_stateElements_10 <= mulContext_delay_17_stateElements_10;
    mulContext_delay_19_isFull <= mulContext_delay_18_isFull;
    mulContext_delay_19_fullRound <= mulContext_delay_18_fullRound;
    mulContext_delay_19_partialRound <= mulContext_delay_18_partialRound;
    mulContext_delay_19_stateSize <= mulContext_delay_18_stateSize;
    mulContext_delay_19_stateID <= mulContext_delay_18_stateID;
    mulContext_delay_19_stateElements_0 <= mulContext_delay_18_stateElements_0;
    mulContext_delay_19_stateElements_1 <= mulContext_delay_18_stateElements_1;
    mulContext_delay_19_stateElements_2 <= mulContext_delay_18_stateElements_2;
    mulContext_delay_19_stateElements_3 <= mulContext_delay_18_stateElements_3;
    mulContext_delay_19_stateElements_4 <= mulContext_delay_18_stateElements_4;
    mulContext_delay_19_stateElements_5 <= mulContext_delay_18_stateElements_5;
    mulContext_delay_19_stateElements_6 <= mulContext_delay_18_stateElements_6;
    mulContext_delay_19_stateElements_7 <= mulContext_delay_18_stateElements_7;
    mulContext_delay_19_stateElements_8 <= mulContext_delay_18_stateElements_8;
    mulContext_delay_19_stateElements_9 <= mulContext_delay_18_stateElements_9;
    mulContext_delay_19_stateElements_10 <= mulContext_delay_18_stateElements_10;
    mulContext_delay_20_isFull <= mulContext_delay_19_isFull;
    mulContext_delay_20_fullRound <= mulContext_delay_19_fullRound;
    mulContext_delay_20_partialRound <= mulContext_delay_19_partialRound;
    mulContext_delay_20_stateSize <= mulContext_delay_19_stateSize;
    mulContext_delay_20_stateID <= mulContext_delay_19_stateID;
    mulContext_delay_20_stateElements_0 <= mulContext_delay_19_stateElements_0;
    mulContext_delay_20_stateElements_1 <= mulContext_delay_19_stateElements_1;
    mulContext_delay_20_stateElements_2 <= mulContext_delay_19_stateElements_2;
    mulContext_delay_20_stateElements_3 <= mulContext_delay_19_stateElements_3;
    mulContext_delay_20_stateElements_4 <= mulContext_delay_19_stateElements_4;
    mulContext_delay_20_stateElements_5 <= mulContext_delay_19_stateElements_5;
    mulContext_delay_20_stateElements_6 <= mulContext_delay_19_stateElements_6;
    mulContext_delay_20_stateElements_7 <= mulContext_delay_19_stateElements_7;
    mulContext_delay_20_stateElements_8 <= mulContext_delay_19_stateElements_8;
    mulContext_delay_20_stateElements_9 <= mulContext_delay_19_stateElements_9;
    mulContext_delay_20_stateElements_10 <= mulContext_delay_19_stateElements_10;
    mulContext_delay_21_isFull <= mulContext_delay_20_isFull;
    mulContext_delay_21_fullRound <= mulContext_delay_20_fullRound;
    mulContext_delay_21_partialRound <= mulContext_delay_20_partialRound;
    mulContext_delay_21_stateSize <= mulContext_delay_20_stateSize;
    mulContext_delay_21_stateID <= mulContext_delay_20_stateID;
    mulContext_delay_21_stateElements_0 <= mulContext_delay_20_stateElements_0;
    mulContext_delay_21_stateElements_1 <= mulContext_delay_20_stateElements_1;
    mulContext_delay_21_stateElements_2 <= mulContext_delay_20_stateElements_2;
    mulContext_delay_21_stateElements_3 <= mulContext_delay_20_stateElements_3;
    mulContext_delay_21_stateElements_4 <= mulContext_delay_20_stateElements_4;
    mulContext_delay_21_stateElements_5 <= mulContext_delay_20_stateElements_5;
    mulContext_delay_21_stateElements_6 <= mulContext_delay_20_stateElements_6;
    mulContext_delay_21_stateElements_7 <= mulContext_delay_20_stateElements_7;
    mulContext_delay_21_stateElements_8 <= mulContext_delay_20_stateElements_8;
    mulContext_delay_21_stateElements_9 <= mulContext_delay_20_stateElements_9;
    mulContext_delay_21_stateElements_10 <= mulContext_delay_20_stateElements_10;
    mulContext_delay_22_isFull <= mulContext_delay_21_isFull;
    mulContext_delay_22_fullRound <= mulContext_delay_21_fullRound;
    mulContext_delay_22_partialRound <= mulContext_delay_21_partialRound;
    mulContext_delay_22_stateSize <= mulContext_delay_21_stateSize;
    mulContext_delay_22_stateID <= mulContext_delay_21_stateID;
    mulContext_delay_22_stateElements_0 <= mulContext_delay_21_stateElements_0;
    mulContext_delay_22_stateElements_1 <= mulContext_delay_21_stateElements_1;
    mulContext_delay_22_stateElements_2 <= mulContext_delay_21_stateElements_2;
    mulContext_delay_22_stateElements_3 <= mulContext_delay_21_stateElements_3;
    mulContext_delay_22_stateElements_4 <= mulContext_delay_21_stateElements_4;
    mulContext_delay_22_stateElements_5 <= mulContext_delay_21_stateElements_5;
    mulContext_delay_22_stateElements_6 <= mulContext_delay_21_stateElements_6;
    mulContext_delay_22_stateElements_7 <= mulContext_delay_21_stateElements_7;
    mulContext_delay_22_stateElements_8 <= mulContext_delay_21_stateElements_8;
    mulContext_delay_22_stateElements_9 <= mulContext_delay_21_stateElements_9;
    mulContext_delay_22_stateElements_10 <= mulContext_delay_21_stateElements_10;
    mulContext_delay_23_isFull <= mulContext_delay_22_isFull;
    mulContext_delay_23_fullRound <= mulContext_delay_22_fullRound;
    mulContext_delay_23_partialRound <= mulContext_delay_22_partialRound;
    mulContext_delay_23_stateSize <= mulContext_delay_22_stateSize;
    mulContext_delay_23_stateID <= mulContext_delay_22_stateID;
    mulContext_delay_23_stateElements_0 <= mulContext_delay_22_stateElements_0;
    mulContext_delay_23_stateElements_1 <= mulContext_delay_22_stateElements_1;
    mulContext_delay_23_stateElements_2 <= mulContext_delay_22_stateElements_2;
    mulContext_delay_23_stateElements_3 <= mulContext_delay_22_stateElements_3;
    mulContext_delay_23_stateElements_4 <= mulContext_delay_22_stateElements_4;
    mulContext_delay_23_stateElements_5 <= mulContext_delay_22_stateElements_5;
    mulContext_delay_23_stateElements_6 <= mulContext_delay_22_stateElements_6;
    mulContext_delay_23_stateElements_7 <= mulContext_delay_22_stateElements_7;
    mulContext_delay_23_stateElements_8 <= mulContext_delay_22_stateElements_8;
    mulContext_delay_23_stateElements_9 <= mulContext_delay_22_stateElements_9;
    mulContext_delay_23_stateElements_10 <= mulContext_delay_22_stateElements_10;
    mulContext_delay_24_isFull <= mulContext_delay_23_isFull;
    mulContext_delay_24_fullRound <= mulContext_delay_23_fullRound;
    mulContext_delay_24_partialRound <= mulContext_delay_23_partialRound;
    mulContext_delay_24_stateSize <= mulContext_delay_23_stateSize;
    mulContext_delay_24_stateID <= mulContext_delay_23_stateID;
    mulContext_delay_24_stateElements_0 <= mulContext_delay_23_stateElements_0;
    mulContext_delay_24_stateElements_1 <= mulContext_delay_23_stateElements_1;
    mulContext_delay_24_stateElements_2 <= mulContext_delay_23_stateElements_2;
    mulContext_delay_24_stateElements_3 <= mulContext_delay_23_stateElements_3;
    mulContext_delay_24_stateElements_4 <= mulContext_delay_23_stateElements_4;
    mulContext_delay_24_stateElements_5 <= mulContext_delay_23_stateElements_5;
    mulContext_delay_24_stateElements_6 <= mulContext_delay_23_stateElements_6;
    mulContext_delay_24_stateElements_7 <= mulContext_delay_23_stateElements_7;
    mulContext_delay_24_stateElements_8 <= mulContext_delay_23_stateElements_8;
    mulContext_delay_24_stateElements_9 <= mulContext_delay_23_stateElements_9;
    mulContext_delay_24_stateElements_10 <= mulContext_delay_23_stateElements_10;
    mulContext_delay_25_isFull <= mulContext_delay_24_isFull;
    mulContext_delay_25_fullRound <= mulContext_delay_24_fullRound;
    mulContext_delay_25_partialRound <= mulContext_delay_24_partialRound;
    mulContext_delay_25_stateSize <= mulContext_delay_24_stateSize;
    mulContext_delay_25_stateID <= mulContext_delay_24_stateID;
    mulContext_delay_25_stateElements_0 <= mulContext_delay_24_stateElements_0;
    mulContext_delay_25_stateElements_1 <= mulContext_delay_24_stateElements_1;
    mulContext_delay_25_stateElements_2 <= mulContext_delay_24_stateElements_2;
    mulContext_delay_25_stateElements_3 <= mulContext_delay_24_stateElements_3;
    mulContext_delay_25_stateElements_4 <= mulContext_delay_24_stateElements_4;
    mulContext_delay_25_stateElements_5 <= mulContext_delay_24_stateElements_5;
    mulContext_delay_25_stateElements_6 <= mulContext_delay_24_stateElements_6;
    mulContext_delay_25_stateElements_7 <= mulContext_delay_24_stateElements_7;
    mulContext_delay_25_stateElements_8 <= mulContext_delay_24_stateElements_8;
    mulContext_delay_25_stateElements_9 <= mulContext_delay_24_stateElements_9;
    mulContext_delay_25_stateElements_10 <= mulContext_delay_24_stateElements_10;
    mulContext_delay_26_isFull <= mulContext_delay_25_isFull;
    mulContext_delay_26_fullRound <= mulContext_delay_25_fullRound;
    mulContext_delay_26_partialRound <= mulContext_delay_25_partialRound;
    mulContext_delay_26_stateSize <= mulContext_delay_25_stateSize;
    mulContext_delay_26_stateID <= mulContext_delay_25_stateID;
    mulContext_delay_26_stateElements_0 <= mulContext_delay_25_stateElements_0;
    mulContext_delay_26_stateElements_1 <= mulContext_delay_25_stateElements_1;
    mulContext_delay_26_stateElements_2 <= mulContext_delay_25_stateElements_2;
    mulContext_delay_26_stateElements_3 <= mulContext_delay_25_stateElements_3;
    mulContext_delay_26_stateElements_4 <= mulContext_delay_25_stateElements_4;
    mulContext_delay_26_stateElements_5 <= mulContext_delay_25_stateElements_5;
    mulContext_delay_26_stateElements_6 <= mulContext_delay_25_stateElements_6;
    mulContext_delay_26_stateElements_7 <= mulContext_delay_25_stateElements_7;
    mulContext_delay_26_stateElements_8 <= mulContext_delay_25_stateElements_8;
    mulContext_delay_26_stateElements_9 <= mulContext_delay_25_stateElements_9;
    mulContext_delay_26_stateElements_10 <= mulContext_delay_25_stateElements_10;
    mulContext_delay_27_isFull <= mulContext_delay_26_isFull;
    mulContext_delay_27_fullRound <= mulContext_delay_26_fullRound;
    mulContext_delay_27_partialRound <= mulContext_delay_26_partialRound;
    mulContext_delay_27_stateSize <= mulContext_delay_26_stateSize;
    mulContext_delay_27_stateID <= mulContext_delay_26_stateID;
    mulContext_delay_27_stateElements_0 <= mulContext_delay_26_stateElements_0;
    mulContext_delay_27_stateElements_1 <= mulContext_delay_26_stateElements_1;
    mulContext_delay_27_stateElements_2 <= mulContext_delay_26_stateElements_2;
    mulContext_delay_27_stateElements_3 <= mulContext_delay_26_stateElements_3;
    mulContext_delay_27_stateElements_4 <= mulContext_delay_26_stateElements_4;
    mulContext_delay_27_stateElements_5 <= mulContext_delay_26_stateElements_5;
    mulContext_delay_27_stateElements_6 <= mulContext_delay_26_stateElements_6;
    mulContext_delay_27_stateElements_7 <= mulContext_delay_26_stateElements_7;
    mulContext_delay_27_stateElements_8 <= mulContext_delay_26_stateElements_8;
    mulContext_delay_27_stateElements_9 <= mulContext_delay_26_stateElements_9;
    mulContext_delay_27_stateElements_10 <= mulContext_delay_26_stateElements_10;
    mulContext_delay_28_isFull <= mulContext_delay_27_isFull;
    mulContext_delay_28_fullRound <= mulContext_delay_27_fullRound;
    mulContext_delay_28_partialRound <= mulContext_delay_27_partialRound;
    mulContext_delay_28_stateSize <= mulContext_delay_27_stateSize;
    mulContext_delay_28_stateID <= mulContext_delay_27_stateID;
    mulContext_delay_28_stateElements_0 <= mulContext_delay_27_stateElements_0;
    mulContext_delay_28_stateElements_1 <= mulContext_delay_27_stateElements_1;
    mulContext_delay_28_stateElements_2 <= mulContext_delay_27_stateElements_2;
    mulContext_delay_28_stateElements_3 <= mulContext_delay_27_stateElements_3;
    mulContext_delay_28_stateElements_4 <= mulContext_delay_27_stateElements_4;
    mulContext_delay_28_stateElements_5 <= mulContext_delay_27_stateElements_5;
    mulContext_delay_28_stateElements_6 <= mulContext_delay_27_stateElements_6;
    mulContext_delay_28_stateElements_7 <= mulContext_delay_27_stateElements_7;
    mulContext_delay_28_stateElements_8 <= mulContext_delay_27_stateElements_8;
    mulContext_delay_28_stateElements_9 <= mulContext_delay_27_stateElements_9;
    mulContext_delay_28_stateElements_10 <= mulContext_delay_27_stateElements_10;
    mulContext_delay_29_isFull <= mulContext_delay_28_isFull;
    mulContext_delay_29_fullRound <= mulContext_delay_28_fullRound;
    mulContext_delay_29_partialRound <= mulContext_delay_28_partialRound;
    mulContext_delay_29_stateSize <= mulContext_delay_28_stateSize;
    mulContext_delay_29_stateID <= mulContext_delay_28_stateID;
    mulContext_delay_29_stateElements_0 <= mulContext_delay_28_stateElements_0;
    mulContext_delay_29_stateElements_1 <= mulContext_delay_28_stateElements_1;
    mulContext_delay_29_stateElements_2 <= mulContext_delay_28_stateElements_2;
    mulContext_delay_29_stateElements_3 <= mulContext_delay_28_stateElements_3;
    mulContext_delay_29_stateElements_4 <= mulContext_delay_28_stateElements_4;
    mulContext_delay_29_stateElements_5 <= mulContext_delay_28_stateElements_5;
    mulContext_delay_29_stateElements_6 <= mulContext_delay_28_stateElements_6;
    mulContext_delay_29_stateElements_7 <= mulContext_delay_28_stateElements_7;
    mulContext_delay_29_stateElements_8 <= mulContext_delay_28_stateElements_8;
    mulContext_delay_29_stateElements_9 <= mulContext_delay_28_stateElements_9;
    mulContext_delay_29_stateElements_10 <= mulContext_delay_28_stateElements_10;
    mulContext_delay_30_isFull <= mulContext_delay_29_isFull;
    mulContext_delay_30_fullRound <= mulContext_delay_29_fullRound;
    mulContext_delay_30_partialRound <= mulContext_delay_29_partialRound;
    mulContext_delay_30_stateSize <= mulContext_delay_29_stateSize;
    mulContext_delay_30_stateID <= mulContext_delay_29_stateID;
    mulContext_delay_30_stateElements_0 <= mulContext_delay_29_stateElements_0;
    mulContext_delay_30_stateElements_1 <= mulContext_delay_29_stateElements_1;
    mulContext_delay_30_stateElements_2 <= mulContext_delay_29_stateElements_2;
    mulContext_delay_30_stateElements_3 <= mulContext_delay_29_stateElements_3;
    mulContext_delay_30_stateElements_4 <= mulContext_delay_29_stateElements_4;
    mulContext_delay_30_stateElements_5 <= mulContext_delay_29_stateElements_5;
    mulContext_delay_30_stateElements_6 <= mulContext_delay_29_stateElements_6;
    mulContext_delay_30_stateElements_7 <= mulContext_delay_29_stateElements_7;
    mulContext_delay_30_stateElements_8 <= mulContext_delay_29_stateElements_8;
    mulContext_delay_30_stateElements_9 <= mulContext_delay_29_stateElements_9;
    mulContext_delay_30_stateElements_10 <= mulContext_delay_29_stateElements_10;
    mulContext_delay_31_isFull <= mulContext_delay_30_isFull;
    mulContext_delay_31_fullRound <= mulContext_delay_30_fullRound;
    mulContext_delay_31_partialRound <= mulContext_delay_30_partialRound;
    mulContext_delay_31_stateSize <= mulContext_delay_30_stateSize;
    mulContext_delay_31_stateID <= mulContext_delay_30_stateID;
    mulContext_delay_31_stateElements_0 <= mulContext_delay_30_stateElements_0;
    mulContext_delay_31_stateElements_1 <= mulContext_delay_30_stateElements_1;
    mulContext_delay_31_stateElements_2 <= mulContext_delay_30_stateElements_2;
    mulContext_delay_31_stateElements_3 <= mulContext_delay_30_stateElements_3;
    mulContext_delay_31_stateElements_4 <= mulContext_delay_30_stateElements_4;
    mulContext_delay_31_stateElements_5 <= mulContext_delay_30_stateElements_5;
    mulContext_delay_31_stateElements_6 <= mulContext_delay_30_stateElements_6;
    mulContext_delay_31_stateElements_7 <= mulContext_delay_30_stateElements_7;
    mulContext_delay_31_stateElements_8 <= mulContext_delay_30_stateElements_8;
    mulContext_delay_31_stateElements_9 <= mulContext_delay_30_stateElements_9;
    mulContext_delay_31_stateElements_10 <= mulContext_delay_30_stateElements_10;
    mulContext_delay_32_isFull <= mulContext_delay_31_isFull;
    mulContext_delay_32_fullRound <= mulContext_delay_31_fullRound;
    mulContext_delay_32_partialRound <= mulContext_delay_31_partialRound;
    mulContext_delay_32_stateSize <= mulContext_delay_31_stateSize;
    mulContext_delay_32_stateID <= mulContext_delay_31_stateID;
    mulContext_delay_32_stateElements_0 <= mulContext_delay_31_stateElements_0;
    mulContext_delay_32_stateElements_1 <= mulContext_delay_31_stateElements_1;
    mulContext_delay_32_stateElements_2 <= mulContext_delay_31_stateElements_2;
    mulContext_delay_32_stateElements_3 <= mulContext_delay_31_stateElements_3;
    mulContext_delay_32_stateElements_4 <= mulContext_delay_31_stateElements_4;
    mulContext_delay_32_stateElements_5 <= mulContext_delay_31_stateElements_5;
    mulContext_delay_32_stateElements_6 <= mulContext_delay_31_stateElements_6;
    mulContext_delay_32_stateElements_7 <= mulContext_delay_31_stateElements_7;
    mulContext_delay_32_stateElements_8 <= mulContext_delay_31_stateElements_8;
    mulContext_delay_32_stateElements_9 <= mulContext_delay_31_stateElements_9;
    mulContext_delay_32_stateElements_10 <= mulContext_delay_31_stateElements_10;
    mulContext_delay_33_isFull <= mulContext_delay_32_isFull;
    mulContext_delay_33_fullRound <= mulContext_delay_32_fullRound;
    mulContext_delay_33_partialRound <= mulContext_delay_32_partialRound;
    mulContext_delay_33_stateSize <= mulContext_delay_32_stateSize;
    mulContext_delay_33_stateID <= mulContext_delay_32_stateID;
    mulContext_delay_33_stateElements_0 <= mulContext_delay_32_stateElements_0;
    mulContext_delay_33_stateElements_1 <= mulContext_delay_32_stateElements_1;
    mulContext_delay_33_stateElements_2 <= mulContext_delay_32_stateElements_2;
    mulContext_delay_33_stateElements_3 <= mulContext_delay_32_stateElements_3;
    mulContext_delay_33_stateElements_4 <= mulContext_delay_32_stateElements_4;
    mulContext_delay_33_stateElements_5 <= mulContext_delay_32_stateElements_5;
    mulContext_delay_33_stateElements_6 <= mulContext_delay_32_stateElements_6;
    mulContext_delay_33_stateElements_7 <= mulContext_delay_32_stateElements_7;
    mulContext_delay_33_stateElements_8 <= mulContext_delay_32_stateElements_8;
    mulContext_delay_33_stateElements_9 <= mulContext_delay_32_stateElements_9;
    mulContext_delay_33_stateElements_10 <= mulContext_delay_32_stateElements_10;
    mulContext_delay_34_isFull <= mulContext_delay_33_isFull;
    mulContext_delay_34_fullRound <= mulContext_delay_33_fullRound;
    mulContext_delay_34_partialRound <= mulContext_delay_33_partialRound;
    mulContext_delay_34_stateSize <= mulContext_delay_33_stateSize;
    mulContext_delay_34_stateID <= mulContext_delay_33_stateID;
    mulContext_delay_34_stateElements_0 <= mulContext_delay_33_stateElements_0;
    mulContext_delay_34_stateElements_1 <= mulContext_delay_33_stateElements_1;
    mulContext_delay_34_stateElements_2 <= mulContext_delay_33_stateElements_2;
    mulContext_delay_34_stateElements_3 <= mulContext_delay_33_stateElements_3;
    mulContext_delay_34_stateElements_4 <= mulContext_delay_33_stateElements_4;
    mulContext_delay_34_stateElements_5 <= mulContext_delay_33_stateElements_5;
    mulContext_delay_34_stateElements_6 <= mulContext_delay_33_stateElements_6;
    mulContext_delay_34_stateElements_7 <= mulContext_delay_33_stateElements_7;
    mulContext_delay_34_stateElements_8 <= mulContext_delay_33_stateElements_8;
    mulContext_delay_34_stateElements_9 <= mulContext_delay_33_stateElements_9;
    mulContext_delay_34_stateElements_10 <= mulContext_delay_33_stateElements_10;
    mulContext_delay_35_isFull <= mulContext_delay_34_isFull;
    mulContext_delay_35_fullRound <= mulContext_delay_34_fullRound;
    mulContext_delay_35_partialRound <= mulContext_delay_34_partialRound;
    mulContext_delay_35_stateSize <= mulContext_delay_34_stateSize;
    mulContext_delay_35_stateID <= mulContext_delay_34_stateID;
    mulContext_delay_35_stateElements_0 <= mulContext_delay_34_stateElements_0;
    mulContext_delay_35_stateElements_1 <= mulContext_delay_34_stateElements_1;
    mulContext_delay_35_stateElements_2 <= mulContext_delay_34_stateElements_2;
    mulContext_delay_35_stateElements_3 <= mulContext_delay_34_stateElements_3;
    mulContext_delay_35_stateElements_4 <= mulContext_delay_34_stateElements_4;
    mulContext_delay_35_stateElements_5 <= mulContext_delay_34_stateElements_5;
    mulContext_delay_35_stateElements_6 <= mulContext_delay_34_stateElements_6;
    mulContext_delay_35_stateElements_7 <= mulContext_delay_34_stateElements_7;
    mulContext_delay_35_stateElements_8 <= mulContext_delay_34_stateElements_8;
    mulContext_delay_35_stateElements_9 <= mulContext_delay_34_stateElements_9;
    mulContext_delay_35_stateElements_10 <= mulContext_delay_34_stateElements_10;
    mulContext_delay_36_isFull <= mulContext_delay_35_isFull;
    mulContext_delay_36_fullRound <= mulContext_delay_35_fullRound;
    mulContext_delay_36_partialRound <= mulContext_delay_35_partialRound;
    mulContext_delay_36_stateSize <= mulContext_delay_35_stateSize;
    mulContext_delay_36_stateID <= mulContext_delay_35_stateID;
    mulContext_delay_36_stateElements_0 <= mulContext_delay_35_stateElements_0;
    mulContext_delay_36_stateElements_1 <= mulContext_delay_35_stateElements_1;
    mulContext_delay_36_stateElements_2 <= mulContext_delay_35_stateElements_2;
    mulContext_delay_36_stateElements_3 <= mulContext_delay_35_stateElements_3;
    mulContext_delay_36_stateElements_4 <= mulContext_delay_35_stateElements_4;
    mulContext_delay_36_stateElements_5 <= mulContext_delay_35_stateElements_5;
    mulContext_delay_36_stateElements_6 <= mulContext_delay_35_stateElements_6;
    mulContext_delay_36_stateElements_7 <= mulContext_delay_35_stateElements_7;
    mulContext_delay_36_stateElements_8 <= mulContext_delay_35_stateElements_8;
    mulContext_delay_36_stateElements_9 <= mulContext_delay_35_stateElements_9;
    mulContext_delay_36_stateElements_10 <= mulContext_delay_35_stateElements_10;
    mulContext_delay_37_isFull <= mulContext_delay_36_isFull;
    mulContext_delay_37_fullRound <= mulContext_delay_36_fullRound;
    mulContext_delay_37_partialRound <= mulContext_delay_36_partialRound;
    mulContext_delay_37_stateSize <= mulContext_delay_36_stateSize;
    mulContext_delay_37_stateID <= mulContext_delay_36_stateID;
    mulContext_delay_37_stateElements_0 <= mulContext_delay_36_stateElements_0;
    mulContext_delay_37_stateElements_1 <= mulContext_delay_36_stateElements_1;
    mulContext_delay_37_stateElements_2 <= mulContext_delay_36_stateElements_2;
    mulContext_delay_37_stateElements_3 <= mulContext_delay_36_stateElements_3;
    mulContext_delay_37_stateElements_4 <= mulContext_delay_36_stateElements_4;
    mulContext_delay_37_stateElements_5 <= mulContext_delay_36_stateElements_5;
    mulContext_delay_37_stateElements_6 <= mulContext_delay_36_stateElements_6;
    mulContext_delay_37_stateElements_7 <= mulContext_delay_36_stateElements_7;
    mulContext_delay_37_stateElements_8 <= mulContext_delay_36_stateElements_8;
    mulContext_delay_37_stateElements_9 <= mulContext_delay_36_stateElements_9;
    mulContext_delay_37_stateElements_10 <= mulContext_delay_36_stateElements_10;
    mulContext_delay_38_isFull <= mulContext_delay_37_isFull;
    mulContext_delay_38_fullRound <= mulContext_delay_37_fullRound;
    mulContext_delay_38_partialRound <= mulContext_delay_37_partialRound;
    mulContext_delay_38_stateSize <= mulContext_delay_37_stateSize;
    mulContext_delay_38_stateID <= mulContext_delay_37_stateID;
    mulContext_delay_38_stateElements_0 <= mulContext_delay_37_stateElements_0;
    mulContext_delay_38_stateElements_1 <= mulContext_delay_37_stateElements_1;
    mulContext_delay_38_stateElements_2 <= mulContext_delay_37_stateElements_2;
    mulContext_delay_38_stateElements_3 <= mulContext_delay_37_stateElements_3;
    mulContext_delay_38_stateElements_4 <= mulContext_delay_37_stateElements_4;
    mulContext_delay_38_stateElements_5 <= mulContext_delay_37_stateElements_5;
    mulContext_delay_38_stateElements_6 <= mulContext_delay_37_stateElements_6;
    mulContext_delay_38_stateElements_7 <= mulContext_delay_37_stateElements_7;
    mulContext_delay_38_stateElements_8 <= mulContext_delay_37_stateElements_8;
    mulContext_delay_38_stateElements_9 <= mulContext_delay_37_stateElements_9;
    mulContext_delay_38_stateElements_10 <= mulContext_delay_37_stateElements_10;
    mulContext_delay_39_isFull <= mulContext_delay_38_isFull;
    mulContext_delay_39_fullRound <= mulContext_delay_38_fullRound;
    mulContext_delay_39_partialRound <= mulContext_delay_38_partialRound;
    mulContext_delay_39_stateSize <= mulContext_delay_38_stateSize;
    mulContext_delay_39_stateID <= mulContext_delay_38_stateID;
    mulContext_delay_39_stateElements_0 <= mulContext_delay_38_stateElements_0;
    mulContext_delay_39_stateElements_1 <= mulContext_delay_38_stateElements_1;
    mulContext_delay_39_stateElements_2 <= mulContext_delay_38_stateElements_2;
    mulContext_delay_39_stateElements_3 <= mulContext_delay_38_stateElements_3;
    mulContext_delay_39_stateElements_4 <= mulContext_delay_38_stateElements_4;
    mulContext_delay_39_stateElements_5 <= mulContext_delay_38_stateElements_5;
    mulContext_delay_39_stateElements_6 <= mulContext_delay_38_stateElements_6;
    mulContext_delay_39_stateElements_7 <= mulContext_delay_38_stateElements_7;
    mulContext_delay_39_stateElements_8 <= mulContext_delay_38_stateElements_8;
    mulContext_delay_39_stateElements_9 <= mulContext_delay_38_stateElements_9;
    mulContext_delay_39_stateElements_10 <= mulContext_delay_38_stateElements_10;
    mulContext_delay_40_isFull <= mulContext_delay_39_isFull;
    mulContext_delay_40_fullRound <= mulContext_delay_39_fullRound;
    mulContext_delay_40_partialRound <= mulContext_delay_39_partialRound;
    mulContext_delay_40_stateSize <= mulContext_delay_39_stateSize;
    mulContext_delay_40_stateID <= mulContext_delay_39_stateID;
    mulContext_delay_40_stateElements_0 <= mulContext_delay_39_stateElements_0;
    mulContext_delay_40_stateElements_1 <= mulContext_delay_39_stateElements_1;
    mulContext_delay_40_stateElements_2 <= mulContext_delay_39_stateElements_2;
    mulContext_delay_40_stateElements_3 <= mulContext_delay_39_stateElements_3;
    mulContext_delay_40_stateElements_4 <= mulContext_delay_39_stateElements_4;
    mulContext_delay_40_stateElements_5 <= mulContext_delay_39_stateElements_5;
    mulContext_delay_40_stateElements_6 <= mulContext_delay_39_stateElements_6;
    mulContext_delay_40_stateElements_7 <= mulContext_delay_39_stateElements_7;
    mulContext_delay_40_stateElements_8 <= mulContext_delay_39_stateElements_8;
    mulContext_delay_40_stateElements_9 <= mulContext_delay_39_stateElements_9;
    mulContext_delay_40_stateElements_10 <= mulContext_delay_39_stateElements_10;
    mulContext_delay_41_isFull <= mulContext_delay_40_isFull;
    mulContext_delay_41_fullRound <= mulContext_delay_40_fullRound;
    mulContext_delay_41_partialRound <= mulContext_delay_40_partialRound;
    mulContext_delay_41_stateSize <= mulContext_delay_40_stateSize;
    mulContext_delay_41_stateID <= mulContext_delay_40_stateID;
    mulContext_delay_41_stateElements_0 <= mulContext_delay_40_stateElements_0;
    mulContext_delay_41_stateElements_1 <= mulContext_delay_40_stateElements_1;
    mulContext_delay_41_stateElements_2 <= mulContext_delay_40_stateElements_2;
    mulContext_delay_41_stateElements_3 <= mulContext_delay_40_stateElements_3;
    mulContext_delay_41_stateElements_4 <= mulContext_delay_40_stateElements_4;
    mulContext_delay_41_stateElements_5 <= mulContext_delay_40_stateElements_5;
    mulContext_delay_41_stateElements_6 <= mulContext_delay_40_stateElements_6;
    mulContext_delay_41_stateElements_7 <= mulContext_delay_40_stateElements_7;
    mulContext_delay_41_stateElements_8 <= mulContext_delay_40_stateElements_8;
    mulContext_delay_41_stateElements_9 <= mulContext_delay_40_stateElements_9;
    mulContext_delay_41_stateElements_10 <= mulContext_delay_40_stateElements_10;
    mulContext_delay_42_isFull <= mulContext_delay_41_isFull;
    mulContext_delay_42_fullRound <= mulContext_delay_41_fullRound;
    mulContext_delay_42_partialRound <= mulContext_delay_41_partialRound;
    mulContext_delay_42_stateSize <= mulContext_delay_41_stateSize;
    mulContext_delay_42_stateID <= mulContext_delay_41_stateID;
    mulContext_delay_42_stateElements_0 <= mulContext_delay_41_stateElements_0;
    mulContext_delay_42_stateElements_1 <= mulContext_delay_41_stateElements_1;
    mulContext_delay_42_stateElements_2 <= mulContext_delay_41_stateElements_2;
    mulContext_delay_42_stateElements_3 <= mulContext_delay_41_stateElements_3;
    mulContext_delay_42_stateElements_4 <= mulContext_delay_41_stateElements_4;
    mulContext_delay_42_stateElements_5 <= mulContext_delay_41_stateElements_5;
    mulContext_delay_42_stateElements_6 <= mulContext_delay_41_stateElements_6;
    mulContext_delay_42_stateElements_7 <= mulContext_delay_41_stateElements_7;
    mulContext_delay_42_stateElements_8 <= mulContext_delay_41_stateElements_8;
    mulContext_delay_42_stateElements_9 <= mulContext_delay_41_stateElements_9;
    mulContext_delay_42_stateElements_10 <= mulContext_delay_41_stateElements_10;
    mulContext_delay_43_isFull <= mulContext_delay_42_isFull;
    mulContext_delay_43_fullRound <= mulContext_delay_42_fullRound;
    mulContext_delay_43_partialRound <= mulContext_delay_42_partialRound;
    mulContext_delay_43_stateSize <= mulContext_delay_42_stateSize;
    mulContext_delay_43_stateID <= mulContext_delay_42_stateID;
    mulContext_delay_43_stateElements_0 <= mulContext_delay_42_stateElements_0;
    mulContext_delay_43_stateElements_1 <= mulContext_delay_42_stateElements_1;
    mulContext_delay_43_stateElements_2 <= mulContext_delay_42_stateElements_2;
    mulContext_delay_43_stateElements_3 <= mulContext_delay_42_stateElements_3;
    mulContext_delay_43_stateElements_4 <= mulContext_delay_42_stateElements_4;
    mulContext_delay_43_stateElements_5 <= mulContext_delay_42_stateElements_5;
    mulContext_delay_43_stateElements_6 <= mulContext_delay_42_stateElements_6;
    mulContext_delay_43_stateElements_7 <= mulContext_delay_42_stateElements_7;
    mulContext_delay_43_stateElements_8 <= mulContext_delay_42_stateElements_8;
    mulContext_delay_43_stateElements_9 <= mulContext_delay_42_stateElements_9;
    mulContext_delay_43_stateElements_10 <= mulContext_delay_42_stateElements_10;
    mulContext_delay_44_isFull <= mulContext_delay_43_isFull;
    mulContext_delay_44_fullRound <= mulContext_delay_43_fullRound;
    mulContext_delay_44_partialRound <= mulContext_delay_43_partialRound;
    mulContext_delay_44_stateSize <= mulContext_delay_43_stateSize;
    mulContext_delay_44_stateID <= mulContext_delay_43_stateID;
    mulContext_delay_44_stateElements_0 <= mulContext_delay_43_stateElements_0;
    mulContext_delay_44_stateElements_1 <= mulContext_delay_43_stateElements_1;
    mulContext_delay_44_stateElements_2 <= mulContext_delay_43_stateElements_2;
    mulContext_delay_44_stateElements_3 <= mulContext_delay_43_stateElements_3;
    mulContext_delay_44_stateElements_4 <= mulContext_delay_43_stateElements_4;
    mulContext_delay_44_stateElements_5 <= mulContext_delay_43_stateElements_5;
    mulContext_delay_44_stateElements_6 <= mulContext_delay_43_stateElements_6;
    mulContext_delay_44_stateElements_7 <= mulContext_delay_43_stateElements_7;
    mulContext_delay_44_stateElements_8 <= mulContext_delay_43_stateElements_8;
    mulContext_delay_44_stateElements_9 <= mulContext_delay_43_stateElements_9;
    mulContext_delay_44_stateElements_10 <= mulContext_delay_43_stateElements_10;
    mulContext_delay_45_isFull <= mulContext_delay_44_isFull;
    mulContext_delay_45_fullRound <= mulContext_delay_44_fullRound;
    mulContext_delay_45_partialRound <= mulContext_delay_44_partialRound;
    mulContext_delay_45_stateSize <= mulContext_delay_44_stateSize;
    mulContext_delay_45_stateID <= mulContext_delay_44_stateID;
    mulContext_delay_45_stateElements_0 <= mulContext_delay_44_stateElements_0;
    mulContext_delay_45_stateElements_1 <= mulContext_delay_44_stateElements_1;
    mulContext_delay_45_stateElements_2 <= mulContext_delay_44_stateElements_2;
    mulContext_delay_45_stateElements_3 <= mulContext_delay_44_stateElements_3;
    mulContext_delay_45_stateElements_4 <= mulContext_delay_44_stateElements_4;
    mulContext_delay_45_stateElements_5 <= mulContext_delay_44_stateElements_5;
    mulContext_delay_45_stateElements_6 <= mulContext_delay_44_stateElements_6;
    mulContext_delay_45_stateElements_7 <= mulContext_delay_44_stateElements_7;
    mulContext_delay_45_stateElements_8 <= mulContext_delay_44_stateElements_8;
    mulContext_delay_45_stateElements_9 <= mulContext_delay_44_stateElements_9;
    mulContext_delay_45_stateElements_10 <= mulContext_delay_44_stateElements_10;
    mulContext_delay_46_isFull <= mulContext_delay_45_isFull;
    mulContext_delay_46_fullRound <= mulContext_delay_45_fullRound;
    mulContext_delay_46_partialRound <= mulContext_delay_45_partialRound;
    mulContext_delay_46_stateSize <= mulContext_delay_45_stateSize;
    mulContext_delay_46_stateID <= mulContext_delay_45_stateID;
    mulContext_delay_46_stateElements_0 <= mulContext_delay_45_stateElements_0;
    mulContext_delay_46_stateElements_1 <= mulContext_delay_45_stateElements_1;
    mulContext_delay_46_stateElements_2 <= mulContext_delay_45_stateElements_2;
    mulContext_delay_46_stateElements_3 <= mulContext_delay_45_stateElements_3;
    mulContext_delay_46_stateElements_4 <= mulContext_delay_45_stateElements_4;
    mulContext_delay_46_stateElements_5 <= mulContext_delay_45_stateElements_5;
    mulContext_delay_46_stateElements_6 <= mulContext_delay_45_stateElements_6;
    mulContext_delay_46_stateElements_7 <= mulContext_delay_45_stateElements_7;
    mulContext_delay_46_stateElements_8 <= mulContext_delay_45_stateElements_8;
    mulContext_delay_46_stateElements_9 <= mulContext_delay_45_stateElements_9;
    mulContext_delay_46_stateElements_10 <= mulContext_delay_45_stateElements_10;
    mulContext_delay_47_isFull <= mulContext_delay_46_isFull;
    mulContext_delay_47_fullRound <= mulContext_delay_46_fullRound;
    mulContext_delay_47_partialRound <= mulContext_delay_46_partialRound;
    mulContext_delay_47_stateSize <= mulContext_delay_46_stateSize;
    mulContext_delay_47_stateID <= mulContext_delay_46_stateID;
    mulContext_delay_47_stateElements_0 <= mulContext_delay_46_stateElements_0;
    mulContext_delay_47_stateElements_1 <= mulContext_delay_46_stateElements_1;
    mulContext_delay_47_stateElements_2 <= mulContext_delay_46_stateElements_2;
    mulContext_delay_47_stateElements_3 <= mulContext_delay_46_stateElements_3;
    mulContext_delay_47_stateElements_4 <= mulContext_delay_46_stateElements_4;
    mulContext_delay_47_stateElements_5 <= mulContext_delay_46_stateElements_5;
    mulContext_delay_47_stateElements_6 <= mulContext_delay_46_stateElements_6;
    mulContext_delay_47_stateElements_7 <= mulContext_delay_46_stateElements_7;
    mulContext_delay_47_stateElements_8 <= mulContext_delay_46_stateElements_8;
    mulContext_delay_47_stateElements_9 <= mulContext_delay_46_stateElements_9;
    mulContext_delay_47_stateElements_10 <= mulContext_delay_46_stateElements_10;
    mulContext_delay_48_isFull <= mulContext_delay_47_isFull;
    mulContext_delay_48_fullRound <= mulContext_delay_47_fullRound;
    mulContext_delay_48_partialRound <= mulContext_delay_47_partialRound;
    mulContext_delay_48_stateSize <= mulContext_delay_47_stateSize;
    mulContext_delay_48_stateID <= mulContext_delay_47_stateID;
    mulContext_delay_48_stateElements_0 <= mulContext_delay_47_stateElements_0;
    mulContext_delay_48_stateElements_1 <= mulContext_delay_47_stateElements_1;
    mulContext_delay_48_stateElements_2 <= mulContext_delay_47_stateElements_2;
    mulContext_delay_48_stateElements_3 <= mulContext_delay_47_stateElements_3;
    mulContext_delay_48_stateElements_4 <= mulContext_delay_47_stateElements_4;
    mulContext_delay_48_stateElements_5 <= mulContext_delay_47_stateElements_5;
    mulContext_delay_48_stateElements_6 <= mulContext_delay_47_stateElements_6;
    mulContext_delay_48_stateElements_7 <= mulContext_delay_47_stateElements_7;
    mulContext_delay_48_stateElements_8 <= mulContext_delay_47_stateElements_8;
    mulContext_delay_48_stateElements_9 <= mulContext_delay_47_stateElements_9;
    mulContext_delay_48_stateElements_10 <= mulContext_delay_47_stateElements_10;
    mulContext_delay_49_isFull <= mulContext_delay_48_isFull;
    mulContext_delay_49_fullRound <= mulContext_delay_48_fullRound;
    mulContext_delay_49_partialRound <= mulContext_delay_48_partialRound;
    mulContext_delay_49_stateSize <= mulContext_delay_48_stateSize;
    mulContext_delay_49_stateID <= mulContext_delay_48_stateID;
    mulContext_delay_49_stateElements_0 <= mulContext_delay_48_stateElements_0;
    mulContext_delay_49_stateElements_1 <= mulContext_delay_48_stateElements_1;
    mulContext_delay_49_stateElements_2 <= mulContext_delay_48_stateElements_2;
    mulContext_delay_49_stateElements_3 <= mulContext_delay_48_stateElements_3;
    mulContext_delay_49_stateElements_4 <= mulContext_delay_48_stateElements_4;
    mulContext_delay_49_stateElements_5 <= mulContext_delay_48_stateElements_5;
    mulContext_delay_49_stateElements_6 <= mulContext_delay_48_stateElements_6;
    mulContext_delay_49_stateElements_7 <= mulContext_delay_48_stateElements_7;
    mulContext_delay_49_stateElements_8 <= mulContext_delay_48_stateElements_8;
    mulContext_delay_49_stateElements_9 <= mulContext_delay_48_stateElements_9;
    mulContext_delay_49_stateElements_10 <= mulContext_delay_48_stateElements_10;
    mulContextDelayed_isFull <= mulContext_delay_49_isFull;
    mulContextDelayed_fullRound <= mulContext_delay_49_fullRound;
    mulContextDelayed_partialRound <= mulContext_delay_49_partialRound;
    mulContextDelayed_stateSize <= mulContext_delay_49_stateSize;
    mulContextDelayed_stateID <= mulContext_delay_49_stateID;
    mulContextDelayed_stateElements_0 <= mulContext_delay_49_stateElements_0;
    mulContextDelayed_stateElements_1 <= mulContext_delay_49_stateElements_1;
    mulContextDelayed_stateElements_2 <= mulContext_delay_49_stateElements_2;
    mulContextDelayed_stateElements_3 <= mulContext_delay_49_stateElements_3;
    mulContextDelayed_stateElements_4 <= mulContext_delay_49_stateElements_4;
    mulContextDelayed_stateElements_5 <= mulContext_delay_49_stateElements_5;
    mulContextDelayed_stateElements_6 <= mulContext_delay_49_stateElements_6;
    mulContextDelayed_stateElements_7 <= mulContext_delay_49_stateElements_7;
    mulContextDelayed_stateElements_8 <= mulContext_delay_49_stateElements_8;
    mulContextDelayed_stateElements_9 <= mulContext_delay_49_stateElements_9;
    mulContextDelayed_stateElements_10 <= mulContext_delay_49_stateElements_10;
    montgomeryMultFlow_15_io_output_payload_res_delay_1 <= montgomeryMultFlow_15_io_output_payload_res;
    montgomeryMultFlow_15_io_output_payload_res_delay_2 <= montgomeryMultFlow_15_io_output_payload_res_delay_1;
    montgomeryMultFlow_15_io_output_payload_res_delay_3 <= montgomeryMultFlow_15_io_output_payload_res_delay_2;
    montgomeryMultFlow_15_io_output_payload_res_delay_4 <= montgomeryMultFlow_15_io_output_payload_res_delay_3;
    montgomeryMultFlow_15_io_output_payload_res_delay_5 <= montgomeryMultFlow_15_io_output_payload_res_delay_4;
    montgomeryMultFlow_15_io_output_payload_res_delay_6 <= montgomeryMultFlow_15_io_output_payload_res_delay_5;
    montgomeryMultFlow_15_io_output_payload_res_delay_7 <= montgomeryMultFlow_15_io_output_payload_res_delay_6;
    montgomeryMultFlow_15_io_output_payload_res_delay_8 <= montgomeryMultFlow_15_io_output_payload_res_delay_7;
    montgomeryMultFlow_15_io_output_payload_res_delay_9 <= montgomeryMultFlow_15_io_output_payload_res_delay_8;
    montgomeryMultFlow_15_io_output_payload_res_delay_10 <= montgomeryMultFlow_15_io_output_payload_res_delay_9;
    montgomeryMultFlow_15_io_output_payload_res_delay_11 <= montgomeryMultFlow_15_io_output_payload_res_delay_10;
    montgomeryMultFlow_15_io_output_payload_res_delay_12 <= montgomeryMultFlow_15_io_output_payload_res_delay_11;
    montgomeryMultFlow_15_io_output_payload_res_delay_13 <= montgomeryMultFlow_15_io_output_payload_res_delay_12;
    montgomeryMultFlow_15_io_output_payload_res_delay_14 <= montgomeryMultFlow_15_io_output_payload_res_delay_13;
    montgomeryMultFlow_15_io_output_payload_res_delay_15 <= montgomeryMultFlow_15_io_output_payload_res_delay_14;
    mulOutput0Delayed <= montgomeryMultFlow_15_io_output_payload_res_delay_15;
    addContext_delay_1_isFull <= addContext_isFull;
    addContext_delay_1_fullRound <= addContext_fullRound;
    addContext_delay_1_partialRound <= addContext_partialRound;
    addContext_delay_1_stateSize <= addContext_stateSize;
    addContext_delay_1_stateID <= addContext_stateID;
    addContext_delay_2_isFull <= addContext_delay_1_isFull;
    addContext_delay_2_fullRound <= addContext_delay_1_fullRound;
    addContext_delay_2_partialRound <= addContext_delay_1_partialRound;
    addContext_delay_2_stateSize <= addContext_delay_1_stateSize;
    addContext_delay_2_stateID <= addContext_delay_1_stateID;
    addContext_delay_3_isFull <= addContext_delay_2_isFull;
    addContext_delay_3_fullRound <= addContext_delay_2_fullRound;
    addContext_delay_3_partialRound <= addContext_delay_2_partialRound;
    addContext_delay_3_stateSize <= addContext_delay_2_stateSize;
    addContext_delay_3_stateID <= addContext_delay_2_stateID;
    addContext_delay_4_isFull <= addContext_delay_3_isFull;
    addContext_delay_4_fullRound <= addContext_delay_3_fullRound;
    addContext_delay_4_partialRound <= addContext_delay_3_partialRound;
    addContext_delay_4_stateSize <= addContext_delay_3_stateSize;
    addContext_delay_4_stateID <= addContext_delay_3_stateID;
    addContext_delay_5_isFull <= addContext_delay_4_isFull;
    addContext_delay_5_fullRound <= addContext_delay_4_fullRound;
    addContext_delay_5_partialRound <= addContext_delay_4_partialRound;
    addContext_delay_5_stateSize <= addContext_delay_4_stateSize;
    addContext_delay_5_stateID <= addContext_delay_4_stateID;
    addContext_delay_6_isFull <= addContext_delay_5_isFull;
    addContext_delay_6_fullRound <= addContext_delay_5_fullRound;
    addContext_delay_6_partialRound <= addContext_delay_5_partialRound;
    addContext_delay_6_stateSize <= addContext_delay_5_stateSize;
    addContext_delay_6_stateID <= addContext_delay_5_stateID;
    addContext_delay_7_isFull <= addContext_delay_6_isFull;
    addContext_delay_7_fullRound <= addContext_delay_6_fullRound;
    addContext_delay_7_partialRound <= addContext_delay_6_partialRound;
    addContext_delay_7_stateSize <= addContext_delay_6_stateSize;
    addContext_delay_7_stateID <= addContext_delay_6_stateID;
    addContext_delay_8_isFull <= addContext_delay_7_isFull;
    addContext_delay_8_fullRound <= addContext_delay_7_fullRound;
    addContext_delay_8_partialRound <= addContext_delay_7_partialRound;
    addContext_delay_8_stateSize <= addContext_delay_7_stateSize;
    addContext_delay_8_stateID <= addContext_delay_7_stateID;
    addContext_delay_9_isFull <= addContext_delay_8_isFull;
    addContext_delay_9_fullRound <= addContext_delay_8_fullRound;
    addContext_delay_9_partialRound <= addContext_delay_8_partialRound;
    addContext_delay_9_stateSize <= addContext_delay_8_stateSize;
    addContext_delay_9_stateID <= addContext_delay_8_stateID;
    addContext_delay_10_isFull <= addContext_delay_9_isFull;
    addContext_delay_10_fullRound <= addContext_delay_9_fullRound;
    addContext_delay_10_partialRound <= addContext_delay_9_partialRound;
    addContext_delay_10_stateSize <= addContext_delay_9_stateSize;
    addContext_delay_10_stateID <= addContext_delay_9_stateID;
    addContext_delay_11_isFull <= addContext_delay_10_isFull;
    addContext_delay_11_fullRound <= addContext_delay_10_fullRound;
    addContext_delay_11_partialRound <= addContext_delay_10_partialRound;
    addContext_delay_11_stateSize <= addContext_delay_10_stateSize;
    addContext_delay_11_stateID <= addContext_delay_10_stateID;
    addContext_delay_12_isFull <= addContext_delay_11_isFull;
    addContext_delay_12_fullRound <= addContext_delay_11_fullRound;
    addContext_delay_12_partialRound <= addContext_delay_11_partialRound;
    addContext_delay_12_stateSize <= addContext_delay_11_stateSize;
    addContext_delay_12_stateID <= addContext_delay_11_stateID;
    addContext_delay_13_isFull <= addContext_delay_12_isFull;
    addContext_delay_13_fullRound <= addContext_delay_12_fullRound;
    addContext_delay_13_partialRound <= addContext_delay_12_partialRound;
    addContext_delay_13_stateSize <= addContext_delay_12_stateSize;
    addContext_delay_13_stateID <= addContext_delay_12_stateID;
    addContext_delay_14_isFull <= addContext_delay_13_isFull;
    addContext_delay_14_fullRound <= addContext_delay_13_fullRound;
    addContext_delay_14_partialRound <= addContext_delay_13_partialRound;
    addContext_delay_14_stateSize <= addContext_delay_13_stateSize;
    addContext_delay_14_stateID <= addContext_delay_13_stateID;
    addContext_delay_15_isFull <= addContext_delay_14_isFull;
    addContext_delay_15_fullRound <= addContext_delay_14_fullRound;
    addContext_delay_15_partialRound <= addContext_delay_14_partialRound;
    addContext_delay_15_stateSize <= addContext_delay_14_stateSize;
    addContext_delay_15_stateID <= addContext_delay_14_stateID;
    addContextDelayed_isFull <= addContext_delay_15_isFull;
    addContextDelayed_fullRound <= addContext_delay_15_fullRound;
    addContextDelayed_partialRound <= addContext_delay_15_partialRound;
    addContextDelayed_stateSize <= addContext_delay_15_stateSize;
    addContextDelayed_stateID <= addContext_delay_15_stateID;
  end


endmodule

module ModularAdderFlow (
  input               io_input_valid,
  input      [254:0]  io_input_payload_op1,
  input      [254:0]  io_input_payload_op2,
  output              io_output_valid,
  output     [254:0]  io_output_payload_res,
  input               clk,
  input               resetn
);

  wire                adderIPFlow_4_io_output_valid;
  wire       [255:0]  adderIPFlow_4_io_output_payload_res;
  wire                adderIPFlow_5_io_output_valid;
  wire       [255:0]  adderIPFlow_5_io_output_payload_res;
  wire       [255:0]  _zz__zz_io_output_payload_res;
  wire                adderInput2_valid;
  wire       [254:0]  adderInput2_payload_op1;
  wire       [254:0]  adderInput2_payload_op2;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_1;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_2;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_3;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_4;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_5;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_6;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_7;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_8;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_9;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_10;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_11;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_12;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_13;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_14;
  reg        [255:0]  adderIPFlow_4_io_output_payload_res_delay_15;
  reg        [255:0]  res1Delayed;
  reg                 _zz_io_output_valid;
  reg        [254:0]  _zz_io_output_payload_res;

  assign _zz__zz_io_output_payload_res = ((adderIPFlow_5_io_output_payload_res[255] || res1Delayed[255]) ? adderIPFlow_5_io_output_payload_res : res1Delayed);
  AdderIPFlow adderIPFlow_4 (
    .io_input_valid           (io_input_valid                              ), //i
    .io_input_payload_op1     (io_input_payload_op1[254:0]                 ), //i
    .io_input_payload_op2     (io_input_payload_op2[254:0]                 ), //i
    .io_output_valid          (adderIPFlow_4_io_output_valid               ), //o
    .io_output_payload_res    (adderIPFlow_4_io_output_payload_res[255:0]  ), //o
    .clk                      (clk                                         ), //i
    .resetn                   (resetn                                      )  //i
  );
  AdderIPFlow adderIPFlow_5 (
    .io_input_valid           (adderInput2_valid                           ), //i
    .io_input_payload_op1     (adderInput2_payload_op1[254:0]              ), //i
    .io_input_payload_op2     (adderInput2_payload_op2[254:0]              ), //i
    .io_output_valid          (adderIPFlow_5_io_output_valid               ), //o
    .io_output_payload_res    (adderIPFlow_5_io_output_payload_res[255:0]  ), //o
    .clk                      (clk                                         ), //i
    .resetn                   (resetn                                      )  //i
  );
  assign adderInput2_valid = adderIPFlow_4_io_output_valid;
  assign adderInput2_payload_op1 = adderIPFlow_4_io_output_payload_res[254:0];
  assign adderInput2_payload_op2 = 255'h0c1258acd66282b7ccc627f7f65e27faac425bfd0001a40100000000ffffffff;
  assign io_output_valid = _zz_io_output_valid;
  assign io_output_payload_res = _zz_io_output_payload_res;
  always @(posedge clk) begin
    adderIPFlow_4_io_output_payload_res_delay_1 <= adderIPFlow_4_io_output_payload_res;
    adderIPFlow_4_io_output_payload_res_delay_2 <= adderIPFlow_4_io_output_payload_res_delay_1;
    adderIPFlow_4_io_output_payload_res_delay_3 <= adderIPFlow_4_io_output_payload_res_delay_2;
    adderIPFlow_4_io_output_payload_res_delay_4 <= adderIPFlow_4_io_output_payload_res_delay_3;
    adderIPFlow_4_io_output_payload_res_delay_5 <= adderIPFlow_4_io_output_payload_res_delay_4;
    adderIPFlow_4_io_output_payload_res_delay_6 <= adderIPFlow_4_io_output_payload_res_delay_5;
    adderIPFlow_4_io_output_payload_res_delay_7 <= adderIPFlow_4_io_output_payload_res_delay_6;
    adderIPFlow_4_io_output_payload_res_delay_8 <= adderIPFlow_4_io_output_payload_res_delay_7;
    adderIPFlow_4_io_output_payload_res_delay_9 <= adderIPFlow_4_io_output_payload_res_delay_8;
    adderIPFlow_4_io_output_payload_res_delay_10 <= adderIPFlow_4_io_output_payload_res_delay_9;
    adderIPFlow_4_io_output_payload_res_delay_11 <= adderIPFlow_4_io_output_payload_res_delay_10;
    adderIPFlow_4_io_output_payload_res_delay_12 <= adderIPFlow_4_io_output_payload_res_delay_11;
    adderIPFlow_4_io_output_payload_res_delay_13 <= adderIPFlow_4_io_output_payload_res_delay_12;
    adderIPFlow_4_io_output_payload_res_delay_14 <= adderIPFlow_4_io_output_payload_res_delay_13;
    adderIPFlow_4_io_output_payload_res_delay_15 <= adderIPFlow_4_io_output_payload_res_delay_14;
    res1Delayed <= adderIPFlow_4_io_output_payload_res_delay_15;
    _zz_io_output_payload_res <= _zz__zz_io_output_payload_res[254:0];
  end

  always @(posedge clk) begin
    if(!resetn) begin
      _zz_io_output_valid <= 1'b0;
    end else begin
      _zz_io_output_valid <= adderIPFlow_5_io_output_valid;
    end
  end


endmodule

module RoundConstantMem (
  input               io_addr_isFull,
  input      [2:0]    io_addr_fullRound,
  input      [5:0]    io_addr_partialRound,
  input      [3:0]    io_addr_stateIndex,
  input      [3:0]    io_addr_stateSize,
  output     [254:0]  io_data
);

  wire       [254:0]  fullRoundConstantMem_4_io_constant;
  wire       [254:0]  fullRoundConstantMem_5_io_constant;
  wire       [254:0]  fullRoundConstantMem_6_io_constant;
  wire       [254:0]  fullRoundConstantMem_7_io_constant;
  wire       [254:0]  partialRoundConstantMem_1_io_constant;
  reg        [254:0]  _zz_fullConstant_2;
  wire       [1:0]    _zz_fullConstant_3;
  wire                select_0;
  wire                select_1;
  wire                select_2;
  wire                select_3;
  wire                _zz_fullConstant;
  wire                _zz_fullConstant_1;
  wire       [254:0]  fullConstant;

  assign _zz_fullConstant_3 = {_zz_fullConstant_1,_zz_fullConstant};
  FullRoundConstantMem fullRoundConstantMem_4 (
    .io_stateIndex    (io_addr_stateIndex[3:0]                    ), //i
    .io_fullRound     (io_addr_fullRound[2:0]                     ), //i
    .io_constant      (fullRoundConstantMem_4_io_constant[254:0]  )  //o
  );
  FullRoundConstantMem_1 fullRoundConstantMem_5 (
    .io_stateIndex    (io_addr_stateIndex[3:0]                    ), //i
    .io_fullRound     (io_addr_fullRound[2:0]                     ), //i
    .io_constant      (fullRoundConstantMem_5_io_constant[254:0]  )  //o
  );
  FullRoundConstantMem_2 fullRoundConstantMem_6 (
    .io_stateIndex    (io_addr_stateIndex[3:0]                    ), //i
    .io_fullRound     (io_addr_fullRound[2:0]                     ), //i
    .io_constant      (fullRoundConstantMem_6_io_constant[254:0]  )  //o
  );
  FullRoundConstantMem_3 fullRoundConstantMem_7 (
    .io_stateIndex    (io_addr_stateIndex[3:0]                    ), //i
    .io_fullRound     (io_addr_fullRound[2:0]                     ), //i
    .io_constant      (fullRoundConstantMem_7_io_constant[254:0]  )  //o
  );
  PartialRoundConstantMem partialRoundConstantMem_1 (
    .io_stateSize       (io_addr_stateSize[3:0]                        ), //i
    .io_partialRound    (io_addr_partialRound[5:0]                     ), //i
    .io_constant        (partialRoundConstantMem_1_io_constant[254:0]  )  //o
  );
  always @(*) begin
    case(_zz_fullConstant_3)
      2'b00 : _zz_fullConstant_2 = fullRoundConstantMem_4_io_constant;
      2'b01 : _zz_fullConstant_2 = fullRoundConstantMem_5_io_constant;
      2'b10 : _zz_fullConstant_2 = fullRoundConstantMem_6_io_constant;
      default : _zz_fullConstant_2 = fullRoundConstantMem_7_io_constant;
    endcase
  end

  assign select_0 = (4'b0011 == io_addr_stateSize);
  assign select_1 = (4'b0101 == io_addr_stateSize);
  assign select_2 = (4'b1001 == io_addr_stateSize);
  assign select_3 = (4'b1100 == io_addr_stateSize);
  assign _zz_fullConstant = (select_1 || select_3);
  assign _zz_fullConstant_1 = (select_2 || select_3);
  assign fullConstant = _zz_fullConstant_2;
  assign io_data = (io_addr_isFull ? fullConstant : partialRoundConstantMem_1_io_constant);

endmodule

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//AdderIPFlow_2 replaced by AdderIPFlow_2

module AdderIPFlow_2 (
  input               io_input_valid,
  input      [254:0]  io_input_payload_op1,
  input      [254:0]  io_input_payload_op2,
  output              io_output_valid,
  output     [255:0]  io_output_payload_res,
  input               clk,
  input               resetn
);

  wire       [255:0]  simAdderIP_48_io_outputS;
  reg                 io_input_valid_delay_1;
  reg                 io_input_valid_delay_2;
  reg                 io_input_valid_delay_3;
  reg                 io_input_valid_delay_4;
  reg                 io_input_valid_delay_5;
  reg                 io_input_valid_delay_6;
  reg                 io_input_valid_delay_7;
  reg                 validDelayed;

  SimAdderIP simAdderIP_48 (
    .io_inputA     (io_input_payload_op1[254:0]      ), //i
    .io_inputB     (io_input_payload_op2[254:0]      ), //i
    .io_outputS    (simAdderIP_48_io_outputS[255:0]  ), //o
    .clk           (clk                              ), //i
    .resetn        (resetn                           )  //i
  );
  assign io_output_valid = validDelayed;
  assign io_output_payload_res = simAdderIP_48_io_outputS;
  always @(posedge clk) begin
    if(!resetn) begin
      io_input_valid_delay_1 <= 1'b0;
      io_input_valid_delay_2 <= 1'b0;
      io_input_valid_delay_3 <= 1'b0;
      io_input_valid_delay_4 <= 1'b0;
      io_input_valid_delay_5 <= 1'b0;
      io_input_valid_delay_6 <= 1'b0;
      io_input_valid_delay_7 <= 1'b0;
      validDelayed <= 1'b0;
    end else begin
      io_input_valid_delay_1 <= io_input_valid;
      io_input_valid_delay_2 <= io_input_valid_delay_1;
      io_input_valid_delay_3 <= io_input_valid_delay_2;
      io_input_valid_delay_4 <= io_input_valid_delay_3;
      io_input_valid_delay_5 <= io_input_valid_delay_4;
      io_input_valid_delay_6 <= io_input_valid_delay_5;
      io_input_valid_delay_7 <= io_input_valid_delay_6;
      validDelayed <= io_input_valid_delay_7;
    end
  end


endmodule

module ShiftMatrix (
  input               io_input_valid,
  input               io_input_payload_isFull,
  input      [2:0]    io_input_payload_fullRound,
  input      [5:0]    io_input_payload_partialRound,
  input      [3:0]    io_input_payload_stateSize,
  input      [7:0]    io_input_payload_stateID,
  input      [254:0]  io_input_payload_stateElements_0,
  input      [254:0]  io_input_payload_stateElements_1,
  input      [254:0]  io_input_payload_stateElements_2,
  input      [254:0]  io_input_payload_stateElements_3,
  input      [254:0]  io_input_payload_stateElements_4,
  input      [254:0]  io_input_payload_stateElements_5,
  input      [254:0]  io_input_payload_stateElements_6,
  input      [254:0]  io_input_payload_stateElements_7,
  input      [254:0]  io_input_payload_stateElements_8,
  input      [254:0]  io_input_payload_stateElements_9,
  input      [254:0]  io_input_payload_stateElements_10,
  input      [254:0]  io_input_payload_stateElements_11,
  output reg          io_output_valid,
  output              io_output_payload_isFull,
  output     [2:0]    io_output_payload_fullRound,
  output     [5:0]    io_output_payload_partialRound,
  output     [3:0]    io_output_payload_stateSize,
  output     [7:0]    io_output_payload_stateID,
  output reg [254:0]  io_output_payload_stateElements_0,
  output reg [254:0]  io_output_payload_stateElements_1,
  output reg [254:0]  io_output_payload_stateElements_2,
  output reg [254:0]  io_output_payload_stateElements_3,
  output reg [254:0]  io_output_payload_stateElements_4,
  output reg [254:0]  io_output_payload_stateElements_5,
  output reg [254:0]  io_output_payload_stateElements_6,
  output reg [254:0]  io_output_payload_stateElements_7,
  output reg [254:0]  io_output_payload_stateElements_8,
  output reg [254:0]  io_output_payload_stateElements_9,
  output reg [254:0]  io_output_payload_stateElements_10,
  output reg [254:0]  io_output_payload_stateElements_11,
  input               clk,
  input               resetn
);
  localparam fsm_enumDef_1_BOOT = 3'd0;
  localparam fsm_enumDef_1_R0R1 = 3'd1;
  localparam fsm_enumDef_1_R1R0 = 3'd2;
  localparam fsm_enumDef_1_T0R1 = 3'd3;
  localparam fsm_enumDef_1_R0T1 = 3'd4;

  wire       [254:0]  bufferVec0_0_io_parallelInput_0;
  wire       [254:0]  bufferVec0_0_io_parallelInput_1;
  wire       [254:0]  bufferVec0_0_io_parallelInput_2;
  wire       [254:0]  bufferVec0_0_io_parallelInput_3;
  wire       [254:0]  bufferVec0_0_io_parallelInput_4;
  wire       [254:0]  bufferVec0_0_io_parallelInput_5;
  wire       [254:0]  bufferVec0_0_io_parallelInput_6;
  wire       [254:0]  bufferVec0_0_io_parallelInput_7;
  wire       [254:0]  bufferVec0_0_io_parallelInput_8;
  wire       [254:0]  bufferVec0_0_io_parallelInput_9;
  wire       [254:0]  bufferVec0_0_io_parallelInput_10;
  wire       [254:0]  bufferVec0_0_io_parallelInput_11;
  wire       [254:0]  bufferVec0_1_io_parallelInput_0;
  wire       [254:0]  bufferVec0_1_io_parallelInput_1;
  wire       [254:0]  bufferVec0_1_io_parallelInput_2;
  wire       [254:0]  bufferVec0_1_io_parallelInput_3;
  wire       [254:0]  bufferVec0_1_io_parallelInput_4;
  wire       [254:0]  bufferVec0_1_io_parallelInput_5;
  wire       [254:0]  bufferVec0_1_io_parallelInput_6;
  wire       [254:0]  bufferVec0_1_io_parallelInput_7;
  wire       [254:0]  bufferVec0_1_io_parallelInput_8;
  wire       [254:0]  bufferVec0_1_io_parallelInput_9;
  wire       [254:0]  bufferVec0_1_io_parallelInput_10;
  wire       [254:0]  bufferVec0_1_io_parallelInput_11;
  wire       [254:0]  bufferVec0_2_io_parallelInput_0;
  wire       [254:0]  bufferVec0_2_io_parallelInput_1;
  wire       [254:0]  bufferVec0_2_io_parallelInput_2;
  wire       [254:0]  bufferVec0_2_io_parallelInput_3;
  wire       [254:0]  bufferVec0_2_io_parallelInput_4;
  wire       [254:0]  bufferVec0_2_io_parallelInput_5;
  wire       [254:0]  bufferVec0_2_io_parallelInput_6;
  wire       [254:0]  bufferVec0_2_io_parallelInput_7;
  wire       [254:0]  bufferVec0_2_io_parallelInput_8;
  wire       [254:0]  bufferVec0_2_io_parallelInput_9;
  wire       [254:0]  bufferVec0_2_io_parallelInput_10;
  wire       [254:0]  bufferVec0_2_io_parallelInput_11;
  wire       [254:0]  bufferVec0_3_io_parallelInput_0;
  wire       [254:0]  bufferVec0_3_io_parallelInput_1;
  wire       [254:0]  bufferVec0_3_io_parallelInput_2;
  wire       [254:0]  bufferVec0_3_io_parallelInput_3;
  wire       [254:0]  bufferVec0_3_io_parallelInput_4;
  wire       [254:0]  bufferVec0_3_io_parallelInput_5;
  wire       [254:0]  bufferVec0_3_io_parallelInput_6;
  wire       [254:0]  bufferVec0_3_io_parallelInput_7;
  wire       [254:0]  bufferVec0_3_io_parallelInput_8;
  wire       [254:0]  bufferVec0_3_io_parallelInput_9;
  wire       [254:0]  bufferVec0_3_io_parallelInput_10;
  wire       [254:0]  bufferVec0_3_io_parallelInput_11;
  wire       [254:0]  bufferVec0_4_io_parallelInput_0;
  wire       [254:0]  bufferVec0_4_io_parallelInput_1;
  wire       [254:0]  bufferVec0_4_io_parallelInput_2;
  wire       [254:0]  bufferVec0_4_io_parallelInput_3;
  wire       [254:0]  bufferVec0_4_io_parallelInput_4;
  wire       [254:0]  bufferVec0_4_io_parallelInput_5;
  wire       [254:0]  bufferVec0_4_io_parallelInput_6;
  wire       [254:0]  bufferVec0_4_io_parallelInput_7;
  wire       [254:0]  bufferVec0_4_io_parallelInput_8;
  wire       [254:0]  bufferVec0_4_io_parallelInput_9;
  wire       [254:0]  bufferVec0_4_io_parallelInput_10;
  wire       [254:0]  bufferVec0_4_io_parallelInput_11;
  wire       [254:0]  bufferVec0_5_io_parallelInput_0;
  wire       [254:0]  bufferVec0_5_io_parallelInput_1;
  wire       [254:0]  bufferVec0_5_io_parallelInput_2;
  wire       [254:0]  bufferVec0_5_io_parallelInput_3;
  wire       [254:0]  bufferVec0_5_io_parallelInput_4;
  wire       [254:0]  bufferVec0_5_io_parallelInput_5;
  wire       [254:0]  bufferVec0_5_io_parallelInput_6;
  wire       [254:0]  bufferVec0_5_io_parallelInput_7;
  wire       [254:0]  bufferVec0_5_io_parallelInput_8;
  wire       [254:0]  bufferVec0_5_io_parallelInput_9;
  wire       [254:0]  bufferVec0_5_io_parallelInput_10;
  wire       [254:0]  bufferVec0_5_io_parallelInput_11;
  wire       [254:0]  bufferVec0_6_io_parallelInput_0;
  wire       [254:0]  bufferVec0_6_io_parallelInput_1;
  wire       [254:0]  bufferVec0_6_io_parallelInput_2;
  wire       [254:0]  bufferVec0_6_io_parallelInput_3;
  wire       [254:0]  bufferVec0_6_io_parallelInput_4;
  wire       [254:0]  bufferVec0_6_io_parallelInput_5;
  wire       [254:0]  bufferVec0_6_io_parallelInput_6;
  wire       [254:0]  bufferVec0_6_io_parallelInput_7;
  wire       [254:0]  bufferVec0_6_io_parallelInput_8;
  wire       [254:0]  bufferVec0_6_io_parallelInput_9;
  wire       [254:0]  bufferVec0_6_io_parallelInput_10;
  wire       [254:0]  bufferVec0_6_io_parallelInput_11;
  wire       [254:0]  bufferVec0_7_io_parallelInput_0;
  wire       [254:0]  bufferVec0_7_io_parallelInput_1;
  wire       [254:0]  bufferVec0_7_io_parallelInput_2;
  wire       [254:0]  bufferVec0_7_io_parallelInput_3;
  wire       [254:0]  bufferVec0_7_io_parallelInput_4;
  wire       [254:0]  bufferVec0_7_io_parallelInput_5;
  wire       [254:0]  bufferVec0_7_io_parallelInput_6;
  wire       [254:0]  bufferVec0_7_io_parallelInput_7;
  wire       [254:0]  bufferVec0_7_io_parallelInput_8;
  wire       [254:0]  bufferVec0_7_io_parallelInput_9;
  wire       [254:0]  bufferVec0_7_io_parallelInput_10;
  wire       [254:0]  bufferVec0_7_io_parallelInput_11;
  wire       [254:0]  bufferVec0_8_io_parallelInput_0;
  wire       [254:0]  bufferVec0_8_io_parallelInput_1;
  wire       [254:0]  bufferVec0_8_io_parallelInput_2;
  wire       [254:0]  bufferVec0_8_io_parallelInput_3;
  wire       [254:0]  bufferVec0_8_io_parallelInput_4;
  wire       [254:0]  bufferVec0_8_io_parallelInput_5;
  wire       [254:0]  bufferVec0_8_io_parallelInput_6;
  wire       [254:0]  bufferVec0_8_io_parallelInput_7;
  wire       [254:0]  bufferVec0_8_io_parallelInput_8;
  wire       [254:0]  bufferVec0_8_io_parallelInput_9;
  wire       [254:0]  bufferVec0_8_io_parallelInput_10;
  wire       [254:0]  bufferVec0_8_io_parallelInput_11;
  wire       [254:0]  bufferVec0_9_io_parallelInput_0;
  wire       [254:0]  bufferVec0_9_io_parallelInput_1;
  wire       [254:0]  bufferVec0_9_io_parallelInput_2;
  wire       [254:0]  bufferVec0_9_io_parallelInput_3;
  wire       [254:0]  bufferVec0_9_io_parallelInput_4;
  wire       [254:0]  bufferVec0_9_io_parallelInput_5;
  wire       [254:0]  bufferVec0_9_io_parallelInput_6;
  wire       [254:0]  bufferVec0_9_io_parallelInput_7;
  wire       [254:0]  bufferVec0_9_io_parallelInput_8;
  wire       [254:0]  bufferVec0_9_io_parallelInput_9;
  wire       [254:0]  bufferVec0_9_io_parallelInput_10;
  wire       [254:0]  bufferVec0_9_io_parallelInput_11;
  wire       [254:0]  bufferVec0_10_io_parallelInput_0;
  wire       [254:0]  bufferVec0_10_io_parallelInput_1;
  wire       [254:0]  bufferVec0_10_io_parallelInput_2;
  wire       [254:0]  bufferVec0_10_io_parallelInput_3;
  wire       [254:0]  bufferVec0_10_io_parallelInput_4;
  wire       [254:0]  bufferVec0_10_io_parallelInput_5;
  wire       [254:0]  bufferVec0_10_io_parallelInput_6;
  wire       [254:0]  bufferVec0_10_io_parallelInput_7;
  wire       [254:0]  bufferVec0_10_io_parallelInput_8;
  wire       [254:0]  bufferVec0_10_io_parallelInput_9;
  wire       [254:0]  bufferVec0_10_io_parallelInput_10;
  wire       [254:0]  bufferVec0_10_io_parallelInput_11;
  wire       [254:0]  bufferVec0_11_io_parallelInput_0;
  wire       [254:0]  bufferVec0_11_io_parallelInput_1;
  wire       [254:0]  bufferVec0_11_io_parallelInput_2;
  wire       [254:0]  bufferVec0_11_io_parallelInput_3;
  wire       [254:0]  bufferVec0_11_io_parallelInput_4;
  wire       [254:0]  bufferVec0_11_io_parallelInput_5;
  wire       [254:0]  bufferVec0_11_io_parallelInput_6;
  wire       [254:0]  bufferVec0_11_io_parallelInput_7;
  wire       [254:0]  bufferVec0_11_io_parallelInput_8;
  wire       [254:0]  bufferVec0_11_io_parallelInput_9;
  wire       [254:0]  bufferVec0_11_io_parallelInput_10;
  wire       [254:0]  bufferVec0_11_io_parallelInput_11;
  wire       [254:0]  bufferVec1_0_io_parallelInput_0;
  wire       [254:0]  bufferVec1_0_io_parallelInput_1;
  wire       [254:0]  bufferVec1_0_io_parallelInput_2;
  wire       [254:0]  bufferVec1_0_io_parallelInput_3;
  wire       [254:0]  bufferVec1_0_io_parallelInput_4;
  wire       [254:0]  bufferVec1_0_io_parallelInput_5;
  wire       [254:0]  bufferVec1_0_io_parallelInput_6;
  wire       [254:0]  bufferVec1_0_io_parallelInput_7;
  wire       [254:0]  bufferVec1_0_io_parallelInput_8;
  wire       [254:0]  bufferVec1_0_io_parallelInput_9;
  wire       [254:0]  bufferVec1_0_io_parallelInput_10;
  wire       [254:0]  bufferVec1_0_io_parallelInput_11;
  wire       [254:0]  bufferVec1_1_io_parallelInput_0;
  wire       [254:0]  bufferVec1_1_io_parallelInput_1;
  wire       [254:0]  bufferVec1_1_io_parallelInput_2;
  wire       [254:0]  bufferVec1_1_io_parallelInput_3;
  wire       [254:0]  bufferVec1_1_io_parallelInput_4;
  wire       [254:0]  bufferVec1_1_io_parallelInput_5;
  wire       [254:0]  bufferVec1_1_io_parallelInput_6;
  wire       [254:0]  bufferVec1_1_io_parallelInput_7;
  wire       [254:0]  bufferVec1_1_io_parallelInput_8;
  wire       [254:0]  bufferVec1_1_io_parallelInput_9;
  wire       [254:0]  bufferVec1_1_io_parallelInput_10;
  wire       [254:0]  bufferVec1_1_io_parallelInput_11;
  wire       [254:0]  bufferVec1_2_io_parallelInput_0;
  wire       [254:0]  bufferVec1_2_io_parallelInput_1;
  wire       [254:0]  bufferVec1_2_io_parallelInput_2;
  wire       [254:0]  bufferVec1_2_io_parallelInput_3;
  wire       [254:0]  bufferVec1_2_io_parallelInput_4;
  wire       [254:0]  bufferVec1_2_io_parallelInput_5;
  wire       [254:0]  bufferVec1_2_io_parallelInput_6;
  wire       [254:0]  bufferVec1_2_io_parallelInput_7;
  wire       [254:0]  bufferVec1_2_io_parallelInput_8;
  wire       [254:0]  bufferVec1_2_io_parallelInput_9;
  wire       [254:0]  bufferVec1_2_io_parallelInput_10;
  wire       [254:0]  bufferVec1_2_io_parallelInput_11;
  wire       [254:0]  bufferVec1_3_io_parallelInput_0;
  wire       [254:0]  bufferVec1_3_io_parallelInput_1;
  wire       [254:0]  bufferVec1_3_io_parallelInput_2;
  wire       [254:0]  bufferVec1_3_io_parallelInput_3;
  wire       [254:0]  bufferVec1_3_io_parallelInput_4;
  wire       [254:0]  bufferVec1_3_io_parallelInput_5;
  wire       [254:0]  bufferVec1_3_io_parallelInput_6;
  wire       [254:0]  bufferVec1_3_io_parallelInput_7;
  wire       [254:0]  bufferVec1_3_io_parallelInput_8;
  wire       [254:0]  bufferVec1_3_io_parallelInput_9;
  wire       [254:0]  bufferVec1_3_io_parallelInput_10;
  wire       [254:0]  bufferVec1_3_io_parallelInput_11;
  wire       [254:0]  bufferVec1_4_io_parallelInput_0;
  wire       [254:0]  bufferVec1_4_io_parallelInput_1;
  wire       [254:0]  bufferVec1_4_io_parallelInput_2;
  wire       [254:0]  bufferVec1_4_io_parallelInput_3;
  wire       [254:0]  bufferVec1_4_io_parallelInput_4;
  wire       [254:0]  bufferVec1_4_io_parallelInput_5;
  wire       [254:0]  bufferVec1_4_io_parallelInput_6;
  wire       [254:0]  bufferVec1_4_io_parallelInput_7;
  wire       [254:0]  bufferVec1_4_io_parallelInput_8;
  wire       [254:0]  bufferVec1_4_io_parallelInput_9;
  wire       [254:0]  bufferVec1_4_io_parallelInput_10;
  wire       [254:0]  bufferVec1_4_io_parallelInput_11;
  wire       [254:0]  bufferVec1_5_io_parallelInput_0;
  wire       [254:0]  bufferVec1_5_io_parallelInput_1;
  wire       [254:0]  bufferVec1_5_io_parallelInput_2;
  wire       [254:0]  bufferVec1_5_io_parallelInput_3;
  wire       [254:0]  bufferVec1_5_io_parallelInput_4;
  wire       [254:0]  bufferVec1_5_io_parallelInput_5;
  wire       [254:0]  bufferVec1_5_io_parallelInput_6;
  wire       [254:0]  bufferVec1_5_io_parallelInput_7;
  wire       [254:0]  bufferVec1_5_io_parallelInput_8;
  wire       [254:0]  bufferVec1_5_io_parallelInput_9;
  wire       [254:0]  bufferVec1_5_io_parallelInput_10;
  wire       [254:0]  bufferVec1_5_io_parallelInput_11;
  wire       [254:0]  bufferVec1_6_io_parallelInput_0;
  wire       [254:0]  bufferVec1_6_io_parallelInput_1;
  wire       [254:0]  bufferVec1_6_io_parallelInput_2;
  wire       [254:0]  bufferVec1_6_io_parallelInput_3;
  wire       [254:0]  bufferVec1_6_io_parallelInput_4;
  wire       [254:0]  bufferVec1_6_io_parallelInput_5;
  wire       [254:0]  bufferVec1_6_io_parallelInput_6;
  wire       [254:0]  bufferVec1_6_io_parallelInput_7;
  wire       [254:0]  bufferVec1_6_io_parallelInput_8;
  wire       [254:0]  bufferVec1_6_io_parallelInput_9;
  wire       [254:0]  bufferVec1_6_io_parallelInput_10;
  wire       [254:0]  bufferVec1_6_io_parallelInput_11;
  wire       [254:0]  bufferVec1_7_io_parallelInput_0;
  wire       [254:0]  bufferVec1_7_io_parallelInput_1;
  wire       [254:0]  bufferVec1_7_io_parallelInput_2;
  wire       [254:0]  bufferVec1_7_io_parallelInput_3;
  wire       [254:0]  bufferVec1_7_io_parallelInput_4;
  wire       [254:0]  bufferVec1_7_io_parallelInput_5;
  wire       [254:0]  bufferVec1_7_io_parallelInput_6;
  wire       [254:0]  bufferVec1_7_io_parallelInput_7;
  wire       [254:0]  bufferVec1_7_io_parallelInput_8;
  wire       [254:0]  bufferVec1_7_io_parallelInput_9;
  wire       [254:0]  bufferVec1_7_io_parallelInput_10;
  wire       [254:0]  bufferVec1_7_io_parallelInput_11;
  wire       [254:0]  bufferVec1_8_io_parallelInput_0;
  wire       [254:0]  bufferVec1_8_io_parallelInput_1;
  wire       [254:0]  bufferVec1_8_io_parallelInput_2;
  wire       [254:0]  bufferVec1_8_io_parallelInput_3;
  wire       [254:0]  bufferVec1_8_io_parallelInput_4;
  wire       [254:0]  bufferVec1_8_io_parallelInput_5;
  wire       [254:0]  bufferVec1_8_io_parallelInput_6;
  wire       [254:0]  bufferVec1_8_io_parallelInput_7;
  wire       [254:0]  bufferVec1_8_io_parallelInput_8;
  wire       [254:0]  bufferVec1_8_io_parallelInput_9;
  wire       [254:0]  bufferVec1_8_io_parallelInput_10;
  wire       [254:0]  bufferVec1_8_io_parallelInput_11;
  wire       [254:0]  bufferVec1_9_io_parallelInput_0;
  wire       [254:0]  bufferVec1_9_io_parallelInput_1;
  wire       [254:0]  bufferVec1_9_io_parallelInput_2;
  wire       [254:0]  bufferVec1_9_io_parallelInput_3;
  wire       [254:0]  bufferVec1_9_io_parallelInput_4;
  wire       [254:0]  bufferVec1_9_io_parallelInput_5;
  wire       [254:0]  bufferVec1_9_io_parallelInput_6;
  wire       [254:0]  bufferVec1_9_io_parallelInput_7;
  wire       [254:0]  bufferVec1_9_io_parallelInput_8;
  wire       [254:0]  bufferVec1_9_io_parallelInput_9;
  wire       [254:0]  bufferVec1_9_io_parallelInput_10;
  wire       [254:0]  bufferVec1_9_io_parallelInput_11;
  wire       [254:0]  bufferVec1_10_io_parallelInput_0;
  wire       [254:0]  bufferVec1_10_io_parallelInput_1;
  wire       [254:0]  bufferVec1_10_io_parallelInput_2;
  wire       [254:0]  bufferVec1_10_io_parallelInput_3;
  wire       [254:0]  bufferVec1_10_io_parallelInput_4;
  wire       [254:0]  bufferVec1_10_io_parallelInput_5;
  wire       [254:0]  bufferVec1_10_io_parallelInput_6;
  wire       [254:0]  bufferVec1_10_io_parallelInput_7;
  wire       [254:0]  bufferVec1_10_io_parallelInput_8;
  wire       [254:0]  bufferVec1_10_io_parallelInput_9;
  wire       [254:0]  bufferVec1_10_io_parallelInput_10;
  wire       [254:0]  bufferVec1_10_io_parallelInput_11;
  wire       [254:0]  bufferVec1_11_io_parallelInput_0;
  wire       [254:0]  bufferVec1_11_io_parallelInput_1;
  wire       [254:0]  bufferVec1_11_io_parallelInput_2;
  wire       [254:0]  bufferVec1_11_io_parallelInput_3;
  wire       [254:0]  bufferVec1_11_io_parallelInput_4;
  wire       [254:0]  bufferVec1_11_io_parallelInput_5;
  wire       [254:0]  bufferVec1_11_io_parallelInput_6;
  wire       [254:0]  bufferVec1_11_io_parallelInput_7;
  wire       [254:0]  bufferVec1_11_io_parallelInput_8;
  wire       [254:0]  bufferVec1_11_io_parallelInput_9;
  wire       [254:0]  bufferVec1_11_io_parallelInput_10;
  wire       [254:0]  bufferVec1_11_io_parallelInput_11;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_0_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_1_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_2_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_3_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_4_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_5_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_6_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_7_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_8_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_9_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_10_io_parallelOutput_11;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_0;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_1;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_2;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_3;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_4;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_5;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_6;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_7;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_8;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_9;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_10;
  wire       [254:0]  bufferVec0_11_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_0_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_1_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_2_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_3_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_4_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_5_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_6_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_7_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_8_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_9_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_10_io_parallelOutput_11;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_0;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_1;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_2;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_3;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_4;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_5;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_6;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_7;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_8;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_9;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_10;
  wire       [254:0]  bufferVec1_11_io_parallelOutput_11;
  wire       [254:0]  _zz__zz_io_parallelInput_0;
  wire       [254:0]  _zz__zz_io_parallelInput_0_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_1_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_1_2;
  wire       [254:0]  _zz__zz_io_parallelInput_0_2;
  wire       [254:0]  _zz__zz_io_parallelInput_0_2_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_3;
  wire       [254:0]  _zz__zz_io_parallelInput_0_3_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_4;
  wire       [254:0]  _zz__zz_io_parallelInput_0_4_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_5;
  wire       [254:0]  _zz__zz_io_parallelInput_0_5_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_6;
  wire       [254:0]  _zz__zz_io_parallelInput_0_6_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_7;
  wire       [254:0]  _zz__zz_io_parallelInput_0_7_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_8;
  wire       [254:0]  _zz__zz_io_parallelInput_0_8_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_9;
  wire       [254:0]  _zz__zz_io_parallelInput_0_9_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_10;
  wire       [254:0]  _zz__zz_io_parallelInput_0_10_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_11;
  wire       [254:0]  _zz__zz_io_parallelInput_0_11_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_12;
  wire       [254:0]  _zz__zz_io_parallelInput_0_12_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_13;
  wire       [254:0]  _zz__zz_io_parallelInput_0_13_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_14;
  wire       [254:0]  _zz__zz_io_parallelInput_0_14_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_15;
  wire       [254:0]  _zz__zz_io_parallelInput_0_15_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_16;
  wire       [254:0]  _zz__zz_io_parallelInput_0_16_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_17;
  wire       [254:0]  _zz__zz_io_parallelInput_0_17_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_18;
  wire       [254:0]  _zz__zz_io_parallelInput_0_18_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_19;
  wire       [254:0]  _zz__zz_io_parallelInput_0_19_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_20;
  wire       [254:0]  _zz__zz_io_parallelInput_0_20_1;
  wire       [254:0]  _zz__zz_io_parallelInput_0_21;
  wire       [254:0]  _zz__zz_io_parallelInput_0_21_1;
  wire       [3:0]    _zz_when_MDSMatrixAdders_l257;
  wire       [3:0]    _zz_when_MDSMatrixAdders_l270;
  wire       [254:0]  _zz__zz_io_output_payload_stateElements_0_1;
  wire       [254:0]  _zz__zz_io_output_payload_stateElements_0_1_1;
  wire       [3:0]    _zz_when_MDSMatrixAdders_l292;
  wire       [3:0]    _zz_when_MDSMatrixAdders_l296;
  wire       [254:0]  _zz__zz_io_output_payload_stateElements_0_2;
  wire       [254:0]  _zz__zz_io_output_payload_stateElements_0_2_1;
  wire       [3:0]    _zz_when_MDSMatrixAdders_l317;
  wire       [3:0]    _zz_when_MDSMatrixAdders_l321;
  reg                 bufferEna0;
  reg                 bufferEna1;
  reg                 bufferInit0;
  reg                 bufferInit1;
  wire       [3059:0] _zz_io_parallelInput_0;
  wire       [3059:0] _zz_io_parallelInput_0_1;
  wire       [3059:0] _zz_io_parallelInput_0_2;
  wire       [3059:0] _zz_io_parallelInput_0_3;
  wire       [3059:0] _zz_io_parallelInput_0_4;
  wire       [3059:0] _zz_io_parallelInput_0_5;
  wire       [3059:0] _zz_io_parallelInput_0_6;
  wire       [3059:0] _zz_io_parallelInput_0_7;
  wire       [3059:0] _zz_io_parallelInput_0_8;
  wire       [3059:0] _zz_io_parallelInput_0_9;
  wire       [3059:0] _zz_io_parallelInput_0_10;
  wire       [3059:0] _zz_io_parallelInput_0_11;
  wire       [3059:0] _zz_io_parallelInput_0_12;
  wire       [3059:0] _zz_io_parallelInput_0_13;
  wire       [3059:0] _zz_io_parallelInput_0_14;
  wire       [3059:0] _zz_io_parallelInput_0_15;
  wire       [3059:0] _zz_io_parallelInput_0_16;
  wire       [3059:0] _zz_io_parallelInput_0_17;
  wire       [3059:0] _zz_io_parallelInput_0_18;
  wire       [3059:0] _zz_io_parallelInput_0_19;
  wire       [3059:0] _zz_io_parallelInput_0_20;
  wire       [3059:0] _zz_io_parallelInput_0_21;
  wire       [3059:0] _zz_io_parallelInput_0_22;
  wire       [3059:0] _zz_io_parallelInput_0_23;
  wire                fsm_wantExit;
  reg                 fsm_wantStart;
  wire                fsm_wantKill;
  reg                 fsm_outContext_isFull;
  reg        [2:0]    fsm_outContext_fullRound;
  reg        [5:0]    fsm_outContext_partialRound;
  reg        [3:0]    fsm_outContext_stateSize;
  reg        [7:0]    fsm_outContext_stateID;
  reg        [3:0]    fsm_inCount;
  reg        [3:0]    fsm_outCount;
  wire       [3059:0] _zz_io_output_payload_stateElements_0;
  reg        [2:0]    fsm_stateReg;
  reg        [2:0]    fsm_stateNext;
  wire                when_MDSMatrixAdders_l257;
  wire                when_MDSMatrixAdders_l270;
  wire       [3059:0] _zz_io_output_payload_stateElements_0_1;
  wire                when_MDSMatrixAdders_l292;
  wire                when_MDSMatrixAdders_l296;
  wire       [3059:0] _zz_io_output_payload_stateElements_0_2;
  wire                when_MDSMatrixAdders_l317;
  wire                when_MDSMatrixAdders_l321;
  wire                when_StateMachine_l222;
  wire                when_StateMachine_l222_1;
  wire                when_StateMachine_l222_2;
  wire                when_StateMachine_l222_3;
  `ifndef SYNTHESIS
  reg [31:0] fsm_stateReg_string;
  reg [31:0] fsm_stateNext_string;
  `endif


  assign _zz_when_MDSMatrixAdders_l257 = (io_input_payload_stateSize - 4'b0001);
  assign _zz_when_MDSMatrixAdders_l270 = (io_input_payload_stateSize - 4'b0001);
  assign _zz_when_MDSMatrixAdders_l292 = (io_input_payload_stateSize - 4'b0001);
  assign _zz_when_MDSMatrixAdders_l296 = (fsm_outContext_stateSize - 4'b0001);
  assign _zz_when_MDSMatrixAdders_l317 = (io_input_payload_stateSize - 4'b0001);
  assign _zz_when_MDSMatrixAdders_l321 = (fsm_outContext_stateSize - 4'b0001);
  assign _zz__zz_io_parallelInput_0 = bufferVec0_1_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_1 = bufferVec0_1_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_1_1 = bufferVec1_1_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_1_2 = bufferVec1_1_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_2 = bufferVec0_2_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_2_1 = bufferVec0_2_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_3 = bufferVec1_2_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_3_1 = bufferVec1_2_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_4 = bufferVec0_3_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_4_1 = bufferVec0_3_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_5 = bufferVec1_3_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_5_1 = bufferVec1_3_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_6 = bufferVec0_4_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_6_1 = bufferVec0_4_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_7 = bufferVec1_4_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_7_1 = bufferVec1_4_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_8 = bufferVec0_5_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_8_1 = bufferVec0_5_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_9 = bufferVec1_5_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_9_1 = bufferVec1_5_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_10 = bufferVec0_6_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_10_1 = bufferVec0_6_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_11 = bufferVec1_6_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_11_1 = bufferVec1_6_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_12 = bufferVec0_7_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_12_1 = bufferVec0_7_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_13 = bufferVec1_7_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_13_1 = bufferVec1_7_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_14 = bufferVec0_8_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_14_1 = bufferVec0_8_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_15 = bufferVec1_8_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_15_1 = bufferVec1_8_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_16 = bufferVec0_9_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_16_1 = bufferVec0_9_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_17 = bufferVec1_9_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_17_1 = bufferVec1_9_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_18 = bufferVec0_10_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_18_1 = bufferVec0_10_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_19 = bufferVec1_10_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_19_1 = bufferVec1_10_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_20 = bufferVec0_11_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_20_1 = bufferVec0_11_io_parallelOutput_0;
  assign _zz__zz_io_parallelInput_0_21 = bufferVec1_11_io_parallelOutput_1;
  assign _zz__zz_io_parallelInput_0_21_1 = bufferVec1_11_io_parallelOutput_0;
  assign _zz__zz_io_output_payload_stateElements_0_1 = bufferVec0_0_io_parallelOutput_1;
  assign _zz__zz_io_output_payload_stateElements_0_1_1 = bufferVec0_0_io_parallelOutput_0;
  assign _zz__zz_io_output_payload_stateElements_0_2 = bufferVec1_0_io_parallelOutput_1;
  assign _zz__zz_io_output_payload_stateElements_0_2_1 = bufferVec1_0_io_parallelOutput_0;
  ShiftRegister bufferVec0_0 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_0[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_0_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_0_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_0_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_0_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_0_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_0_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_0_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_0_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_0_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_0_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_0_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_0_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_0_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_0_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_0_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_0_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_0_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_0_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_0_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_0_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_0_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_0_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_0_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_0_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_1 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_1[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_1_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_1_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_1_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_1_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_1_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_1_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_1_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_1_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_1_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_1_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_1_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_1_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_1_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_1_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_1_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_1_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_1_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_1_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_1_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_1_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_1_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_1_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_1_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_1_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_2 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_2[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_2_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_2_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_2_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_2_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_2_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_2_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_2_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_2_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_2_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_2_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_2_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_2_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_2_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_2_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_2_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_2_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_2_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_2_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_2_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_2_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_2_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_2_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_2_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_2_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_3 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_3[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_3_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_3_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_3_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_3_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_3_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_3_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_3_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_3_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_3_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_3_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_3_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_3_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_3_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_3_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_3_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_3_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_3_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_3_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_3_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_3_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_3_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_3_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_3_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_3_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_4 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_4[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_4_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_4_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_4_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_4_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_4_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_4_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_4_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_4_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_4_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_4_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_4_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_4_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_4_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_4_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_4_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_4_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_4_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_4_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_4_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_4_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_4_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_4_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_4_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_4_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_5 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_5[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_5_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_5_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_5_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_5_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_5_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_5_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_5_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_5_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_5_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_5_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_5_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_5_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_5_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_5_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_5_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_5_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_5_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_5_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_5_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_5_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_5_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_5_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_5_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_5_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_6 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_6[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_6_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_6_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_6_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_6_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_6_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_6_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_6_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_6_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_6_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_6_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_6_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_6_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_6_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_6_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_6_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_6_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_6_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_6_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_6_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_6_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_6_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_6_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_6_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_6_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_7 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_7[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_7_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_7_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_7_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_7_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_7_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_7_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_7_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_7_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_7_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_7_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_7_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_7_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_7_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_7_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_7_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_7_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_7_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_7_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_7_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_7_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_7_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_7_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_7_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_7_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_8 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_8[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_8_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_8_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_8_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_8_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_8_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_8_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_8_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_8_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_8_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_8_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_8_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_8_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_8_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_8_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_8_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_8_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_8_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_8_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_8_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_8_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_8_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_8_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_8_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_8_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_9 (
    .io_ena                  (bufferEna0                                ), //i
    .io_init                 (bufferInit0                               ), //i
    .io_serialInput          (io_input_payload_stateElements_9[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_9_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_9_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_9_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_9_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_9_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_9_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_9_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_9_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_9_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_9_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_9_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_9_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_9_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_9_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_9_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_9_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_9_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_9_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_9_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_9_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_9_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_9_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_9_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_9_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec0_10 (
    .io_ena                  (bufferEna0                                 ), //i
    .io_init                 (bufferInit0                                ), //i
    .io_serialInput          (io_input_payload_stateElements_10[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_10_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_10_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_10_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_10_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_10_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_10_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_10_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_10_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_10_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_10_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_10_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_10_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_10_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_10_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_10_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_10_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_10_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_10_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_10_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_10_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_10_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_10_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_10_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_10_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                        ), //i
    .resetn                  (resetn                                     )  //i
  );
  ShiftRegister bufferVec0_11 (
    .io_ena                  (bufferEna0                                 ), //i
    .io_init                 (bufferInit0                                ), //i
    .io_serialInput          (io_input_payload_stateElements_11[254:0]   ), //i
    .io_parallelInput_0      (bufferVec0_11_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec0_11_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec0_11_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec0_11_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec0_11_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec0_11_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec0_11_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec0_11_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec0_11_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec0_11_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec0_11_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec0_11_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec0_11_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec0_11_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec0_11_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec0_11_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec0_11_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec0_11_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec0_11_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec0_11_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec0_11_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec0_11_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec0_11_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec0_11_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                        ), //i
    .resetn                  (resetn                                     )  //i
  );
  ShiftRegister bufferVec1_0 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_0[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_0_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_0_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_0_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_0_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_0_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_0_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_0_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_0_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_0_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_0_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_0_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_0_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_0_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_0_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_0_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_0_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_0_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_0_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_0_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_0_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_0_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_0_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_0_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_0_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_1 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_1[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_1_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_1_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_1_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_1_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_1_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_1_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_1_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_1_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_1_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_1_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_1_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_1_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_1_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_1_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_1_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_1_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_1_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_1_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_1_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_1_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_1_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_1_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_1_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_1_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_2 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_2[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_2_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_2_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_2_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_2_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_2_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_2_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_2_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_2_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_2_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_2_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_2_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_2_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_2_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_2_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_2_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_2_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_2_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_2_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_2_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_2_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_2_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_2_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_2_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_2_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_3 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_3[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_3_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_3_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_3_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_3_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_3_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_3_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_3_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_3_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_3_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_3_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_3_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_3_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_3_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_3_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_3_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_3_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_3_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_3_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_3_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_3_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_3_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_3_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_3_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_3_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_4 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_4[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_4_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_4_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_4_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_4_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_4_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_4_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_4_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_4_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_4_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_4_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_4_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_4_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_4_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_4_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_4_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_4_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_4_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_4_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_4_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_4_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_4_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_4_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_4_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_4_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_5 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_5[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_5_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_5_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_5_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_5_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_5_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_5_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_5_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_5_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_5_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_5_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_5_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_5_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_5_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_5_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_5_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_5_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_5_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_5_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_5_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_5_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_5_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_5_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_5_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_5_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_6 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_6[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_6_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_6_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_6_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_6_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_6_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_6_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_6_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_6_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_6_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_6_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_6_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_6_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_6_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_6_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_6_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_6_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_6_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_6_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_6_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_6_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_6_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_6_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_6_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_6_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_7 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_7[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_7_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_7_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_7_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_7_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_7_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_7_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_7_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_7_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_7_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_7_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_7_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_7_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_7_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_7_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_7_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_7_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_7_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_7_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_7_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_7_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_7_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_7_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_7_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_7_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_8 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_8[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_8_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_8_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_8_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_8_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_8_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_8_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_8_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_8_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_8_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_8_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_8_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_8_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_8_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_8_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_8_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_8_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_8_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_8_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_8_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_8_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_8_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_8_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_8_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_8_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_9 (
    .io_ena                  (bufferEna1                                ), //i
    .io_init                 (bufferInit1                               ), //i
    .io_serialInput          (io_input_payload_stateElements_9[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_9_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_9_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_9_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_9_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_9_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_9_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_9_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_9_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_9_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_9_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_9_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_9_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_9_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_9_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_9_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_9_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_9_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_9_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_9_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_9_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_9_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_9_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_9_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_9_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                       ), //i
    .resetn                  (resetn                                    )  //i
  );
  ShiftRegister bufferVec1_10 (
    .io_ena                  (bufferEna1                                 ), //i
    .io_init                 (bufferInit1                                ), //i
    .io_serialInput          (io_input_payload_stateElements_10[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_10_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_10_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_10_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_10_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_10_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_10_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_10_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_10_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_10_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_10_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_10_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_10_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_10_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_10_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_10_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_10_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_10_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_10_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_10_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_10_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_10_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_10_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_10_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_10_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                        ), //i
    .resetn                  (resetn                                     )  //i
  );
  ShiftRegister bufferVec1_11 (
    .io_ena                  (bufferEna1                                 ), //i
    .io_init                 (bufferInit1                                ), //i
    .io_serialInput          (io_input_payload_stateElements_11[254:0]   ), //i
    .io_parallelInput_0      (bufferVec1_11_io_parallelInput_0[254:0]    ), //i
    .io_parallelInput_1      (bufferVec1_11_io_parallelInput_1[254:0]    ), //i
    .io_parallelInput_2      (bufferVec1_11_io_parallelInput_2[254:0]    ), //i
    .io_parallelInput_3      (bufferVec1_11_io_parallelInput_3[254:0]    ), //i
    .io_parallelInput_4      (bufferVec1_11_io_parallelInput_4[254:0]    ), //i
    .io_parallelInput_5      (bufferVec1_11_io_parallelInput_5[254:0]    ), //i
    .io_parallelInput_6      (bufferVec1_11_io_parallelInput_6[254:0]    ), //i
    .io_parallelInput_7      (bufferVec1_11_io_parallelInput_7[254:0]    ), //i
    .io_parallelInput_8      (bufferVec1_11_io_parallelInput_8[254:0]    ), //i
    .io_parallelInput_9      (bufferVec1_11_io_parallelInput_9[254:0]    ), //i
    .io_parallelInput_10     (bufferVec1_11_io_parallelInput_10[254:0]   ), //i
    .io_parallelInput_11     (bufferVec1_11_io_parallelInput_11[254:0]   ), //i
    .io_parallelOutput_0     (bufferVec1_11_io_parallelOutput_0[254:0]   ), //o
    .io_parallelOutput_1     (bufferVec1_11_io_parallelOutput_1[254:0]   ), //o
    .io_parallelOutput_2     (bufferVec1_11_io_parallelOutput_2[254:0]   ), //o
    .io_parallelOutput_3     (bufferVec1_11_io_parallelOutput_3[254:0]   ), //o
    .io_parallelOutput_4     (bufferVec1_11_io_parallelOutput_4[254:0]   ), //o
    .io_parallelOutput_5     (bufferVec1_11_io_parallelOutput_5[254:0]   ), //o
    .io_parallelOutput_6     (bufferVec1_11_io_parallelOutput_6[254:0]   ), //o
    .io_parallelOutput_7     (bufferVec1_11_io_parallelOutput_7[254:0]   ), //o
    .io_parallelOutput_8     (bufferVec1_11_io_parallelOutput_8[254:0]   ), //o
    .io_parallelOutput_9     (bufferVec1_11_io_parallelOutput_9[254:0]   ), //o
    .io_parallelOutput_10    (bufferVec1_11_io_parallelOutput_10[254:0]  ), //o
    .io_parallelOutput_11    (bufferVec1_11_io_parallelOutput_11[254:0]  ), //o
    .clk                     (clk                                        ), //i
    .resetn                  (resetn                                     )  //i
  );
  `ifndef SYNTHESIS
  always @(*) begin
    case(fsm_stateReg)
      fsm_enumDef_1_BOOT : fsm_stateReg_string = "BOOT";
      fsm_enumDef_1_R0R1 : fsm_stateReg_string = "R0R1";
      fsm_enumDef_1_R1R0 : fsm_stateReg_string = "R1R0";
      fsm_enumDef_1_T0R1 : fsm_stateReg_string = "T0R1";
      fsm_enumDef_1_R0T1 : fsm_stateReg_string = "R0T1";
      default : fsm_stateReg_string = "????";
    endcase
  end
  always @(*) begin
    case(fsm_stateNext)
      fsm_enumDef_1_BOOT : fsm_stateNext_string = "BOOT";
      fsm_enumDef_1_R0R1 : fsm_stateNext_string = "R0R1";
      fsm_enumDef_1_R1R0 : fsm_stateNext_string = "R1R0";
      fsm_enumDef_1_T0R1 : fsm_stateNext_string = "T0R1";
      fsm_enumDef_1_R0T1 : fsm_stateNext_string = "R0T1";
      default : fsm_stateNext_string = "????";
    endcase
  end
  `endif

  assign _zz_io_parallelInput_0 = {bufferVec0_1_io_parallelOutput_11,{bufferVec0_1_io_parallelOutput_10,{bufferVec0_1_io_parallelOutput_9,{bufferVec0_1_io_parallelOutput_8,{bufferVec0_1_io_parallelOutput_7,{bufferVec0_1_io_parallelOutput_6,{bufferVec0_1_io_parallelOutput_5,{bufferVec0_1_io_parallelOutput_4,{bufferVec0_1_io_parallelOutput_3,{bufferVec0_1_io_parallelOutput_2,{_zz__zz_io_parallelInput_0,_zz__zz_io_parallelInput_0_1}}}}}}}}}}};
  assign bufferVec0_0_io_parallelInput_0 = _zz_io_parallelInput_0[254 : 0];
  assign bufferVec0_0_io_parallelInput_1 = _zz_io_parallelInput_0[509 : 255];
  assign bufferVec0_0_io_parallelInput_2 = _zz_io_parallelInput_0[764 : 510];
  assign bufferVec0_0_io_parallelInput_3 = _zz_io_parallelInput_0[1019 : 765];
  assign bufferVec0_0_io_parallelInput_4 = _zz_io_parallelInput_0[1274 : 1020];
  assign bufferVec0_0_io_parallelInput_5 = _zz_io_parallelInput_0[1529 : 1275];
  assign bufferVec0_0_io_parallelInput_6 = _zz_io_parallelInput_0[1784 : 1530];
  assign bufferVec0_0_io_parallelInput_7 = _zz_io_parallelInput_0[2039 : 1785];
  assign bufferVec0_0_io_parallelInput_8 = _zz_io_parallelInput_0[2294 : 2040];
  assign bufferVec0_0_io_parallelInput_9 = _zz_io_parallelInput_0[2549 : 2295];
  assign bufferVec0_0_io_parallelInput_10 = _zz_io_parallelInput_0[2804 : 2550];
  assign bufferVec0_0_io_parallelInput_11 = _zz_io_parallelInput_0[3059 : 2805];
  assign _zz_io_parallelInput_0_1 = {bufferVec1_1_io_parallelOutput_11,{bufferVec1_1_io_parallelOutput_10,{bufferVec1_1_io_parallelOutput_9,{bufferVec1_1_io_parallelOutput_8,{bufferVec1_1_io_parallelOutput_7,{bufferVec1_1_io_parallelOutput_6,{bufferVec1_1_io_parallelOutput_5,{bufferVec1_1_io_parallelOutput_4,{bufferVec1_1_io_parallelOutput_3,{bufferVec1_1_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_1_1,_zz__zz_io_parallelInput_0_1_2}}}}}}}}}}};
  assign bufferVec1_0_io_parallelInput_0 = _zz_io_parallelInput_0_1[254 : 0];
  assign bufferVec1_0_io_parallelInput_1 = _zz_io_parallelInput_0_1[509 : 255];
  assign bufferVec1_0_io_parallelInput_2 = _zz_io_parallelInput_0_1[764 : 510];
  assign bufferVec1_0_io_parallelInput_3 = _zz_io_parallelInput_0_1[1019 : 765];
  assign bufferVec1_0_io_parallelInput_4 = _zz_io_parallelInput_0_1[1274 : 1020];
  assign bufferVec1_0_io_parallelInput_5 = _zz_io_parallelInput_0_1[1529 : 1275];
  assign bufferVec1_0_io_parallelInput_6 = _zz_io_parallelInput_0_1[1784 : 1530];
  assign bufferVec1_0_io_parallelInput_7 = _zz_io_parallelInput_0_1[2039 : 1785];
  assign bufferVec1_0_io_parallelInput_8 = _zz_io_parallelInput_0_1[2294 : 2040];
  assign bufferVec1_0_io_parallelInput_9 = _zz_io_parallelInput_0_1[2549 : 2295];
  assign bufferVec1_0_io_parallelInput_10 = _zz_io_parallelInput_0_1[2804 : 2550];
  assign bufferVec1_0_io_parallelInput_11 = _zz_io_parallelInput_0_1[3059 : 2805];
  assign _zz_io_parallelInput_0_2 = {bufferVec0_2_io_parallelOutput_11,{bufferVec0_2_io_parallelOutput_10,{bufferVec0_2_io_parallelOutput_9,{bufferVec0_2_io_parallelOutput_8,{bufferVec0_2_io_parallelOutput_7,{bufferVec0_2_io_parallelOutput_6,{bufferVec0_2_io_parallelOutput_5,{bufferVec0_2_io_parallelOutput_4,{bufferVec0_2_io_parallelOutput_3,{bufferVec0_2_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_2,_zz__zz_io_parallelInput_0_2_1}}}}}}}}}}};
  assign bufferVec0_1_io_parallelInput_0 = _zz_io_parallelInput_0_2[254 : 0];
  assign bufferVec0_1_io_parallelInput_1 = _zz_io_parallelInput_0_2[509 : 255];
  assign bufferVec0_1_io_parallelInput_2 = _zz_io_parallelInput_0_2[764 : 510];
  assign bufferVec0_1_io_parallelInput_3 = _zz_io_parallelInput_0_2[1019 : 765];
  assign bufferVec0_1_io_parallelInput_4 = _zz_io_parallelInput_0_2[1274 : 1020];
  assign bufferVec0_1_io_parallelInput_5 = _zz_io_parallelInput_0_2[1529 : 1275];
  assign bufferVec0_1_io_parallelInput_6 = _zz_io_parallelInput_0_2[1784 : 1530];
  assign bufferVec0_1_io_parallelInput_7 = _zz_io_parallelInput_0_2[2039 : 1785];
  assign bufferVec0_1_io_parallelInput_8 = _zz_io_parallelInput_0_2[2294 : 2040];
  assign bufferVec0_1_io_parallelInput_9 = _zz_io_parallelInput_0_2[2549 : 2295];
  assign bufferVec0_1_io_parallelInput_10 = _zz_io_parallelInput_0_2[2804 : 2550];
  assign bufferVec0_1_io_parallelInput_11 = _zz_io_parallelInput_0_2[3059 : 2805];
  assign _zz_io_parallelInput_0_3 = {bufferVec1_2_io_parallelOutput_11,{bufferVec1_2_io_parallelOutput_10,{bufferVec1_2_io_parallelOutput_9,{bufferVec1_2_io_parallelOutput_8,{bufferVec1_2_io_parallelOutput_7,{bufferVec1_2_io_parallelOutput_6,{bufferVec1_2_io_parallelOutput_5,{bufferVec1_2_io_parallelOutput_4,{bufferVec1_2_io_parallelOutput_3,{bufferVec1_2_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_3,_zz__zz_io_parallelInput_0_3_1}}}}}}}}}}};
  assign bufferVec1_1_io_parallelInput_0 = _zz_io_parallelInput_0_3[254 : 0];
  assign bufferVec1_1_io_parallelInput_1 = _zz_io_parallelInput_0_3[509 : 255];
  assign bufferVec1_1_io_parallelInput_2 = _zz_io_parallelInput_0_3[764 : 510];
  assign bufferVec1_1_io_parallelInput_3 = _zz_io_parallelInput_0_3[1019 : 765];
  assign bufferVec1_1_io_parallelInput_4 = _zz_io_parallelInput_0_3[1274 : 1020];
  assign bufferVec1_1_io_parallelInput_5 = _zz_io_parallelInput_0_3[1529 : 1275];
  assign bufferVec1_1_io_parallelInput_6 = _zz_io_parallelInput_0_3[1784 : 1530];
  assign bufferVec1_1_io_parallelInput_7 = _zz_io_parallelInput_0_3[2039 : 1785];
  assign bufferVec1_1_io_parallelInput_8 = _zz_io_parallelInput_0_3[2294 : 2040];
  assign bufferVec1_1_io_parallelInput_9 = _zz_io_parallelInput_0_3[2549 : 2295];
  assign bufferVec1_1_io_parallelInput_10 = _zz_io_parallelInput_0_3[2804 : 2550];
  assign bufferVec1_1_io_parallelInput_11 = _zz_io_parallelInput_0_3[3059 : 2805];
  assign _zz_io_parallelInput_0_4 = {bufferVec0_3_io_parallelOutput_11,{bufferVec0_3_io_parallelOutput_10,{bufferVec0_3_io_parallelOutput_9,{bufferVec0_3_io_parallelOutput_8,{bufferVec0_3_io_parallelOutput_7,{bufferVec0_3_io_parallelOutput_6,{bufferVec0_3_io_parallelOutput_5,{bufferVec0_3_io_parallelOutput_4,{bufferVec0_3_io_parallelOutput_3,{bufferVec0_3_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_4,_zz__zz_io_parallelInput_0_4_1}}}}}}}}}}};
  assign bufferVec0_2_io_parallelInput_0 = _zz_io_parallelInput_0_4[254 : 0];
  assign bufferVec0_2_io_parallelInput_1 = _zz_io_parallelInput_0_4[509 : 255];
  assign bufferVec0_2_io_parallelInput_2 = _zz_io_parallelInput_0_4[764 : 510];
  assign bufferVec0_2_io_parallelInput_3 = _zz_io_parallelInput_0_4[1019 : 765];
  assign bufferVec0_2_io_parallelInput_4 = _zz_io_parallelInput_0_4[1274 : 1020];
  assign bufferVec0_2_io_parallelInput_5 = _zz_io_parallelInput_0_4[1529 : 1275];
  assign bufferVec0_2_io_parallelInput_6 = _zz_io_parallelInput_0_4[1784 : 1530];
  assign bufferVec0_2_io_parallelInput_7 = _zz_io_parallelInput_0_4[2039 : 1785];
  assign bufferVec0_2_io_parallelInput_8 = _zz_io_parallelInput_0_4[2294 : 2040];
  assign bufferVec0_2_io_parallelInput_9 = _zz_io_parallelInput_0_4[2549 : 2295];
  assign bufferVec0_2_io_parallelInput_10 = _zz_io_parallelInput_0_4[2804 : 2550];
  assign bufferVec0_2_io_parallelInput_11 = _zz_io_parallelInput_0_4[3059 : 2805];
  assign _zz_io_parallelInput_0_5 = {bufferVec1_3_io_parallelOutput_11,{bufferVec1_3_io_parallelOutput_10,{bufferVec1_3_io_parallelOutput_9,{bufferVec1_3_io_parallelOutput_8,{bufferVec1_3_io_parallelOutput_7,{bufferVec1_3_io_parallelOutput_6,{bufferVec1_3_io_parallelOutput_5,{bufferVec1_3_io_parallelOutput_4,{bufferVec1_3_io_parallelOutput_3,{bufferVec1_3_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_5,_zz__zz_io_parallelInput_0_5_1}}}}}}}}}}};
  assign bufferVec1_2_io_parallelInput_0 = _zz_io_parallelInput_0_5[254 : 0];
  assign bufferVec1_2_io_parallelInput_1 = _zz_io_parallelInput_0_5[509 : 255];
  assign bufferVec1_2_io_parallelInput_2 = _zz_io_parallelInput_0_5[764 : 510];
  assign bufferVec1_2_io_parallelInput_3 = _zz_io_parallelInput_0_5[1019 : 765];
  assign bufferVec1_2_io_parallelInput_4 = _zz_io_parallelInput_0_5[1274 : 1020];
  assign bufferVec1_2_io_parallelInput_5 = _zz_io_parallelInput_0_5[1529 : 1275];
  assign bufferVec1_2_io_parallelInput_6 = _zz_io_parallelInput_0_5[1784 : 1530];
  assign bufferVec1_2_io_parallelInput_7 = _zz_io_parallelInput_0_5[2039 : 1785];
  assign bufferVec1_2_io_parallelInput_8 = _zz_io_parallelInput_0_5[2294 : 2040];
  assign bufferVec1_2_io_parallelInput_9 = _zz_io_parallelInput_0_5[2549 : 2295];
  assign bufferVec1_2_io_parallelInput_10 = _zz_io_parallelInput_0_5[2804 : 2550];
  assign bufferVec1_2_io_parallelInput_11 = _zz_io_parallelInput_0_5[3059 : 2805];
  assign _zz_io_parallelInput_0_6 = {bufferVec0_4_io_parallelOutput_11,{bufferVec0_4_io_parallelOutput_10,{bufferVec0_4_io_parallelOutput_9,{bufferVec0_4_io_parallelOutput_8,{bufferVec0_4_io_parallelOutput_7,{bufferVec0_4_io_parallelOutput_6,{bufferVec0_4_io_parallelOutput_5,{bufferVec0_4_io_parallelOutput_4,{bufferVec0_4_io_parallelOutput_3,{bufferVec0_4_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_6,_zz__zz_io_parallelInput_0_6_1}}}}}}}}}}};
  assign bufferVec0_3_io_parallelInput_0 = _zz_io_parallelInput_0_6[254 : 0];
  assign bufferVec0_3_io_parallelInput_1 = _zz_io_parallelInput_0_6[509 : 255];
  assign bufferVec0_3_io_parallelInput_2 = _zz_io_parallelInput_0_6[764 : 510];
  assign bufferVec0_3_io_parallelInput_3 = _zz_io_parallelInput_0_6[1019 : 765];
  assign bufferVec0_3_io_parallelInput_4 = _zz_io_parallelInput_0_6[1274 : 1020];
  assign bufferVec0_3_io_parallelInput_5 = _zz_io_parallelInput_0_6[1529 : 1275];
  assign bufferVec0_3_io_parallelInput_6 = _zz_io_parallelInput_0_6[1784 : 1530];
  assign bufferVec0_3_io_parallelInput_7 = _zz_io_parallelInput_0_6[2039 : 1785];
  assign bufferVec0_3_io_parallelInput_8 = _zz_io_parallelInput_0_6[2294 : 2040];
  assign bufferVec0_3_io_parallelInput_9 = _zz_io_parallelInput_0_6[2549 : 2295];
  assign bufferVec0_3_io_parallelInput_10 = _zz_io_parallelInput_0_6[2804 : 2550];
  assign bufferVec0_3_io_parallelInput_11 = _zz_io_parallelInput_0_6[3059 : 2805];
  assign _zz_io_parallelInput_0_7 = {bufferVec1_4_io_parallelOutput_11,{bufferVec1_4_io_parallelOutput_10,{bufferVec1_4_io_parallelOutput_9,{bufferVec1_4_io_parallelOutput_8,{bufferVec1_4_io_parallelOutput_7,{bufferVec1_4_io_parallelOutput_6,{bufferVec1_4_io_parallelOutput_5,{bufferVec1_4_io_parallelOutput_4,{bufferVec1_4_io_parallelOutput_3,{bufferVec1_4_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_7,_zz__zz_io_parallelInput_0_7_1}}}}}}}}}}};
  assign bufferVec1_3_io_parallelInput_0 = _zz_io_parallelInput_0_7[254 : 0];
  assign bufferVec1_3_io_parallelInput_1 = _zz_io_parallelInput_0_7[509 : 255];
  assign bufferVec1_3_io_parallelInput_2 = _zz_io_parallelInput_0_7[764 : 510];
  assign bufferVec1_3_io_parallelInput_3 = _zz_io_parallelInput_0_7[1019 : 765];
  assign bufferVec1_3_io_parallelInput_4 = _zz_io_parallelInput_0_7[1274 : 1020];
  assign bufferVec1_3_io_parallelInput_5 = _zz_io_parallelInput_0_7[1529 : 1275];
  assign bufferVec1_3_io_parallelInput_6 = _zz_io_parallelInput_0_7[1784 : 1530];
  assign bufferVec1_3_io_parallelInput_7 = _zz_io_parallelInput_0_7[2039 : 1785];
  assign bufferVec1_3_io_parallelInput_8 = _zz_io_parallelInput_0_7[2294 : 2040];
  assign bufferVec1_3_io_parallelInput_9 = _zz_io_parallelInput_0_7[2549 : 2295];
  assign bufferVec1_3_io_parallelInput_10 = _zz_io_parallelInput_0_7[2804 : 2550];
  assign bufferVec1_3_io_parallelInput_11 = _zz_io_parallelInput_0_7[3059 : 2805];
  assign _zz_io_parallelInput_0_8 = {bufferVec0_5_io_parallelOutput_11,{bufferVec0_5_io_parallelOutput_10,{bufferVec0_5_io_parallelOutput_9,{bufferVec0_5_io_parallelOutput_8,{bufferVec0_5_io_parallelOutput_7,{bufferVec0_5_io_parallelOutput_6,{bufferVec0_5_io_parallelOutput_5,{bufferVec0_5_io_parallelOutput_4,{bufferVec0_5_io_parallelOutput_3,{bufferVec0_5_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_8,_zz__zz_io_parallelInput_0_8_1}}}}}}}}}}};
  assign bufferVec0_4_io_parallelInput_0 = _zz_io_parallelInput_0_8[254 : 0];
  assign bufferVec0_4_io_parallelInput_1 = _zz_io_parallelInput_0_8[509 : 255];
  assign bufferVec0_4_io_parallelInput_2 = _zz_io_parallelInput_0_8[764 : 510];
  assign bufferVec0_4_io_parallelInput_3 = _zz_io_parallelInput_0_8[1019 : 765];
  assign bufferVec0_4_io_parallelInput_4 = _zz_io_parallelInput_0_8[1274 : 1020];
  assign bufferVec0_4_io_parallelInput_5 = _zz_io_parallelInput_0_8[1529 : 1275];
  assign bufferVec0_4_io_parallelInput_6 = _zz_io_parallelInput_0_8[1784 : 1530];
  assign bufferVec0_4_io_parallelInput_7 = _zz_io_parallelInput_0_8[2039 : 1785];
  assign bufferVec0_4_io_parallelInput_8 = _zz_io_parallelInput_0_8[2294 : 2040];
  assign bufferVec0_4_io_parallelInput_9 = _zz_io_parallelInput_0_8[2549 : 2295];
  assign bufferVec0_4_io_parallelInput_10 = _zz_io_parallelInput_0_8[2804 : 2550];
  assign bufferVec0_4_io_parallelInput_11 = _zz_io_parallelInput_0_8[3059 : 2805];
  assign _zz_io_parallelInput_0_9 = {bufferVec1_5_io_parallelOutput_11,{bufferVec1_5_io_parallelOutput_10,{bufferVec1_5_io_parallelOutput_9,{bufferVec1_5_io_parallelOutput_8,{bufferVec1_5_io_parallelOutput_7,{bufferVec1_5_io_parallelOutput_6,{bufferVec1_5_io_parallelOutput_5,{bufferVec1_5_io_parallelOutput_4,{bufferVec1_5_io_parallelOutput_3,{bufferVec1_5_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_9,_zz__zz_io_parallelInput_0_9_1}}}}}}}}}}};
  assign bufferVec1_4_io_parallelInput_0 = _zz_io_parallelInput_0_9[254 : 0];
  assign bufferVec1_4_io_parallelInput_1 = _zz_io_parallelInput_0_9[509 : 255];
  assign bufferVec1_4_io_parallelInput_2 = _zz_io_parallelInput_0_9[764 : 510];
  assign bufferVec1_4_io_parallelInput_3 = _zz_io_parallelInput_0_9[1019 : 765];
  assign bufferVec1_4_io_parallelInput_4 = _zz_io_parallelInput_0_9[1274 : 1020];
  assign bufferVec1_4_io_parallelInput_5 = _zz_io_parallelInput_0_9[1529 : 1275];
  assign bufferVec1_4_io_parallelInput_6 = _zz_io_parallelInput_0_9[1784 : 1530];
  assign bufferVec1_4_io_parallelInput_7 = _zz_io_parallelInput_0_9[2039 : 1785];
  assign bufferVec1_4_io_parallelInput_8 = _zz_io_parallelInput_0_9[2294 : 2040];
  assign bufferVec1_4_io_parallelInput_9 = _zz_io_parallelInput_0_9[2549 : 2295];
  assign bufferVec1_4_io_parallelInput_10 = _zz_io_parallelInput_0_9[2804 : 2550];
  assign bufferVec1_4_io_parallelInput_11 = _zz_io_parallelInput_0_9[3059 : 2805];
  assign _zz_io_parallelInput_0_10 = {bufferVec0_6_io_parallelOutput_11,{bufferVec0_6_io_parallelOutput_10,{bufferVec0_6_io_parallelOutput_9,{bufferVec0_6_io_parallelOutput_8,{bufferVec0_6_io_parallelOutput_7,{bufferVec0_6_io_parallelOutput_6,{bufferVec0_6_io_parallelOutput_5,{bufferVec0_6_io_parallelOutput_4,{bufferVec0_6_io_parallelOutput_3,{bufferVec0_6_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_10,_zz__zz_io_parallelInput_0_10_1}}}}}}}}}}};
  assign bufferVec0_5_io_parallelInput_0 = _zz_io_parallelInput_0_10[254 : 0];
  assign bufferVec0_5_io_parallelInput_1 = _zz_io_parallelInput_0_10[509 : 255];
  assign bufferVec0_5_io_parallelInput_2 = _zz_io_parallelInput_0_10[764 : 510];
  assign bufferVec0_5_io_parallelInput_3 = _zz_io_parallelInput_0_10[1019 : 765];
  assign bufferVec0_5_io_parallelInput_4 = _zz_io_parallelInput_0_10[1274 : 1020];
  assign bufferVec0_5_io_parallelInput_5 = _zz_io_parallelInput_0_10[1529 : 1275];
  assign bufferVec0_5_io_parallelInput_6 = _zz_io_parallelInput_0_10[1784 : 1530];
  assign bufferVec0_5_io_parallelInput_7 = _zz_io_parallelInput_0_10[2039 : 1785];
  assign bufferVec0_5_io_parallelInput_8 = _zz_io_parallelInput_0_10[2294 : 2040];
  assign bufferVec0_5_io_parallelInput_9 = _zz_io_parallelInput_0_10[2549 : 2295];
  assign bufferVec0_5_io_parallelInput_10 = _zz_io_parallelInput_0_10[2804 : 2550];
  assign bufferVec0_5_io_parallelInput_11 = _zz_io_parallelInput_0_10[3059 : 2805];
  assign _zz_io_parallelInput_0_11 = {bufferVec1_6_io_parallelOutput_11,{bufferVec1_6_io_parallelOutput_10,{bufferVec1_6_io_parallelOutput_9,{bufferVec1_6_io_parallelOutput_8,{bufferVec1_6_io_parallelOutput_7,{bufferVec1_6_io_parallelOutput_6,{bufferVec1_6_io_parallelOutput_5,{bufferVec1_6_io_parallelOutput_4,{bufferVec1_6_io_parallelOutput_3,{bufferVec1_6_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_11,_zz__zz_io_parallelInput_0_11_1}}}}}}}}}}};
  assign bufferVec1_5_io_parallelInput_0 = _zz_io_parallelInput_0_11[254 : 0];
  assign bufferVec1_5_io_parallelInput_1 = _zz_io_parallelInput_0_11[509 : 255];
  assign bufferVec1_5_io_parallelInput_2 = _zz_io_parallelInput_0_11[764 : 510];
  assign bufferVec1_5_io_parallelInput_3 = _zz_io_parallelInput_0_11[1019 : 765];
  assign bufferVec1_5_io_parallelInput_4 = _zz_io_parallelInput_0_11[1274 : 1020];
  assign bufferVec1_5_io_parallelInput_5 = _zz_io_parallelInput_0_11[1529 : 1275];
  assign bufferVec1_5_io_parallelInput_6 = _zz_io_parallelInput_0_11[1784 : 1530];
  assign bufferVec1_5_io_parallelInput_7 = _zz_io_parallelInput_0_11[2039 : 1785];
  assign bufferVec1_5_io_parallelInput_8 = _zz_io_parallelInput_0_11[2294 : 2040];
  assign bufferVec1_5_io_parallelInput_9 = _zz_io_parallelInput_0_11[2549 : 2295];
  assign bufferVec1_5_io_parallelInput_10 = _zz_io_parallelInput_0_11[2804 : 2550];
  assign bufferVec1_5_io_parallelInput_11 = _zz_io_parallelInput_0_11[3059 : 2805];
  assign _zz_io_parallelInput_0_12 = {bufferVec0_7_io_parallelOutput_11,{bufferVec0_7_io_parallelOutput_10,{bufferVec0_7_io_parallelOutput_9,{bufferVec0_7_io_parallelOutput_8,{bufferVec0_7_io_parallelOutput_7,{bufferVec0_7_io_parallelOutput_6,{bufferVec0_7_io_parallelOutput_5,{bufferVec0_7_io_parallelOutput_4,{bufferVec0_7_io_parallelOutput_3,{bufferVec0_7_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_12,_zz__zz_io_parallelInput_0_12_1}}}}}}}}}}};
  assign bufferVec0_6_io_parallelInput_0 = _zz_io_parallelInput_0_12[254 : 0];
  assign bufferVec0_6_io_parallelInput_1 = _zz_io_parallelInput_0_12[509 : 255];
  assign bufferVec0_6_io_parallelInput_2 = _zz_io_parallelInput_0_12[764 : 510];
  assign bufferVec0_6_io_parallelInput_3 = _zz_io_parallelInput_0_12[1019 : 765];
  assign bufferVec0_6_io_parallelInput_4 = _zz_io_parallelInput_0_12[1274 : 1020];
  assign bufferVec0_6_io_parallelInput_5 = _zz_io_parallelInput_0_12[1529 : 1275];
  assign bufferVec0_6_io_parallelInput_6 = _zz_io_parallelInput_0_12[1784 : 1530];
  assign bufferVec0_6_io_parallelInput_7 = _zz_io_parallelInput_0_12[2039 : 1785];
  assign bufferVec0_6_io_parallelInput_8 = _zz_io_parallelInput_0_12[2294 : 2040];
  assign bufferVec0_6_io_parallelInput_9 = _zz_io_parallelInput_0_12[2549 : 2295];
  assign bufferVec0_6_io_parallelInput_10 = _zz_io_parallelInput_0_12[2804 : 2550];
  assign bufferVec0_6_io_parallelInput_11 = _zz_io_parallelInput_0_12[3059 : 2805];
  assign _zz_io_parallelInput_0_13 = {bufferVec1_7_io_parallelOutput_11,{bufferVec1_7_io_parallelOutput_10,{bufferVec1_7_io_parallelOutput_9,{bufferVec1_7_io_parallelOutput_8,{bufferVec1_7_io_parallelOutput_7,{bufferVec1_7_io_parallelOutput_6,{bufferVec1_7_io_parallelOutput_5,{bufferVec1_7_io_parallelOutput_4,{bufferVec1_7_io_parallelOutput_3,{bufferVec1_7_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_13,_zz__zz_io_parallelInput_0_13_1}}}}}}}}}}};
  assign bufferVec1_6_io_parallelInput_0 = _zz_io_parallelInput_0_13[254 : 0];
  assign bufferVec1_6_io_parallelInput_1 = _zz_io_parallelInput_0_13[509 : 255];
  assign bufferVec1_6_io_parallelInput_2 = _zz_io_parallelInput_0_13[764 : 510];
  assign bufferVec1_6_io_parallelInput_3 = _zz_io_parallelInput_0_13[1019 : 765];
  assign bufferVec1_6_io_parallelInput_4 = _zz_io_parallelInput_0_13[1274 : 1020];
  assign bufferVec1_6_io_parallelInput_5 = _zz_io_parallelInput_0_13[1529 : 1275];
  assign bufferVec1_6_io_parallelInput_6 = _zz_io_parallelInput_0_13[1784 : 1530];
  assign bufferVec1_6_io_parallelInput_7 = _zz_io_parallelInput_0_13[2039 : 1785];
  assign bufferVec1_6_io_parallelInput_8 = _zz_io_parallelInput_0_13[2294 : 2040];
  assign bufferVec1_6_io_parallelInput_9 = _zz_io_parallelInput_0_13[2549 : 2295];
  assign bufferVec1_6_io_parallelInput_10 = _zz_io_parallelInput_0_13[2804 : 2550];
  assign bufferVec1_6_io_parallelInput_11 = _zz_io_parallelInput_0_13[3059 : 2805];
  assign _zz_io_parallelInput_0_14 = {bufferVec0_8_io_parallelOutput_11,{bufferVec0_8_io_parallelOutput_10,{bufferVec0_8_io_parallelOutput_9,{bufferVec0_8_io_parallelOutput_8,{bufferVec0_8_io_parallelOutput_7,{bufferVec0_8_io_parallelOutput_6,{bufferVec0_8_io_parallelOutput_5,{bufferVec0_8_io_parallelOutput_4,{bufferVec0_8_io_parallelOutput_3,{bufferVec0_8_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_14,_zz__zz_io_parallelInput_0_14_1}}}}}}}}}}};
  assign bufferVec0_7_io_parallelInput_0 = _zz_io_parallelInput_0_14[254 : 0];
  assign bufferVec0_7_io_parallelInput_1 = _zz_io_parallelInput_0_14[509 : 255];
  assign bufferVec0_7_io_parallelInput_2 = _zz_io_parallelInput_0_14[764 : 510];
  assign bufferVec0_7_io_parallelInput_3 = _zz_io_parallelInput_0_14[1019 : 765];
  assign bufferVec0_7_io_parallelInput_4 = _zz_io_parallelInput_0_14[1274 : 1020];
  assign bufferVec0_7_io_parallelInput_5 = _zz_io_parallelInput_0_14[1529 : 1275];
  assign bufferVec0_7_io_parallelInput_6 = _zz_io_parallelInput_0_14[1784 : 1530];
  assign bufferVec0_7_io_parallelInput_7 = _zz_io_parallelInput_0_14[2039 : 1785];
  assign bufferVec0_7_io_parallelInput_8 = _zz_io_parallelInput_0_14[2294 : 2040];
  assign bufferVec0_7_io_parallelInput_9 = _zz_io_parallelInput_0_14[2549 : 2295];
  assign bufferVec0_7_io_parallelInput_10 = _zz_io_parallelInput_0_14[2804 : 2550];
  assign bufferVec0_7_io_parallelInput_11 = _zz_io_parallelInput_0_14[3059 : 2805];
  assign _zz_io_parallelInput_0_15 = {bufferVec1_8_io_parallelOutput_11,{bufferVec1_8_io_parallelOutput_10,{bufferVec1_8_io_parallelOutput_9,{bufferVec1_8_io_parallelOutput_8,{bufferVec1_8_io_parallelOutput_7,{bufferVec1_8_io_parallelOutput_6,{bufferVec1_8_io_parallelOutput_5,{bufferVec1_8_io_parallelOutput_4,{bufferVec1_8_io_parallelOutput_3,{bufferVec1_8_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_15,_zz__zz_io_parallelInput_0_15_1}}}}}}}}}}};
  assign bufferVec1_7_io_parallelInput_0 = _zz_io_parallelInput_0_15[254 : 0];
  assign bufferVec1_7_io_parallelInput_1 = _zz_io_parallelInput_0_15[509 : 255];
  assign bufferVec1_7_io_parallelInput_2 = _zz_io_parallelInput_0_15[764 : 510];
  assign bufferVec1_7_io_parallelInput_3 = _zz_io_parallelInput_0_15[1019 : 765];
  assign bufferVec1_7_io_parallelInput_4 = _zz_io_parallelInput_0_15[1274 : 1020];
  assign bufferVec1_7_io_parallelInput_5 = _zz_io_parallelInput_0_15[1529 : 1275];
  assign bufferVec1_7_io_parallelInput_6 = _zz_io_parallelInput_0_15[1784 : 1530];
  assign bufferVec1_7_io_parallelInput_7 = _zz_io_parallelInput_0_15[2039 : 1785];
  assign bufferVec1_7_io_parallelInput_8 = _zz_io_parallelInput_0_15[2294 : 2040];
  assign bufferVec1_7_io_parallelInput_9 = _zz_io_parallelInput_0_15[2549 : 2295];
  assign bufferVec1_7_io_parallelInput_10 = _zz_io_parallelInput_0_15[2804 : 2550];
  assign bufferVec1_7_io_parallelInput_11 = _zz_io_parallelInput_0_15[3059 : 2805];
  assign _zz_io_parallelInput_0_16 = {bufferVec0_9_io_parallelOutput_11,{bufferVec0_9_io_parallelOutput_10,{bufferVec0_9_io_parallelOutput_9,{bufferVec0_9_io_parallelOutput_8,{bufferVec0_9_io_parallelOutput_7,{bufferVec0_9_io_parallelOutput_6,{bufferVec0_9_io_parallelOutput_5,{bufferVec0_9_io_parallelOutput_4,{bufferVec0_9_io_parallelOutput_3,{bufferVec0_9_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_16,_zz__zz_io_parallelInput_0_16_1}}}}}}}}}}};
  assign bufferVec0_8_io_parallelInput_0 = _zz_io_parallelInput_0_16[254 : 0];
  assign bufferVec0_8_io_parallelInput_1 = _zz_io_parallelInput_0_16[509 : 255];
  assign bufferVec0_8_io_parallelInput_2 = _zz_io_parallelInput_0_16[764 : 510];
  assign bufferVec0_8_io_parallelInput_3 = _zz_io_parallelInput_0_16[1019 : 765];
  assign bufferVec0_8_io_parallelInput_4 = _zz_io_parallelInput_0_16[1274 : 1020];
  assign bufferVec0_8_io_parallelInput_5 = _zz_io_parallelInput_0_16[1529 : 1275];
  assign bufferVec0_8_io_parallelInput_6 = _zz_io_parallelInput_0_16[1784 : 1530];
  assign bufferVec0_8_io_parallelInput_7 = _zz_io_parallelInput_0_16[2039 : 1785];
  assign bufferVec0_8_io_parallelInput_8 = _zz_io_parallelInput_0_16[2294 : 2040];
  assign bufferVec0_8_io_parallelInput_9 = _zz_io_parallelInput_0_16[2549 : 2295];
  assign bufferVec0_8_io_parallelInput_10 = _zz_io_parallelInput_0_16[2804 : 2550];
  assign bufferVec0_8_io_parallelInput_11 = _zz_io_parallelInput_0_16[3059 : 2805];
  assign _zz_io_parallelInput_0_17 = {bufferVec1_9_io_parallelOutput_11,{bufferVec1_9_io_parallelOutput_10,{bufferVec1_9_io_parallelOutput_9,{bufferVec1_9_io_parallelOutput_8,{bufferVec1_9_io_parallelOutput_7,{bufferVec1_9_io_parallelOutput_6,{bufferVec1_9_io_parallelOutput_5,{bufferVec1_9_io_parallelOutput_4,{bufferVec1_9_io_parallelOutput_3,{bufferVec1_9_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_17,_zz__zz_io_parallelInput_0_17_1}}}}}}}}}}};
  assign bufferVec1_8_io_parallelInput_0 = _zz_io_parallelInput_0_17[254 : 0];
  assign bufferVec1_8_io_parallelInput_1 = _zz_io_parallelInput_0_17[509 : 255];
  assign bufferVec1_8_io_parallelInput_2 = _zz_io_parallelInput_0_17[764 : 510];
  assign bufferVec1_8_io_parallelInput_3 = _zz_io_parallelInput_0_17[1019 : 765];
  assign bufferVec1_8_io_parallelInput_4 = _zz_io_parallelInput_0_17[1274 : 1020];
  assign bufferVec1_8_io_parallelInput_5 = _zz_io_parallelInput_0_17[1529 : 1275];
  assign bufferVec1_8_io_parallelInput_6 = _zz_io_parallelInput_0_17[1784 : 1530];
  assign bufferVec1_8_io_parallelInput_7 = _zz_io_parallelInput_0_17[2039 : 1785];
  assign bufferVec1_8_io_parallelInput_8 = _zz_io_parallelInput_0_17[2294 : 2040];
  assign bufferVec1_8_io_parallelInput_9 = _zz_io_parallelInput_0_17[2549 : 2295];
  assign bufferVec1_8_io_parallelInput_10 = _zz_io_parallelInput_0_17[2804 : 2550];
  assign bufferVec1_8_io_parallelInput_11 = _zz_io_parallelInput_0_17[3059 : 2805];
  assign _zz_io_parallelInput_0_18 = {bufferVec0_10_io_parallelOutput_11,{bufferVec0_10_io_parallelOutput_10,{bufferVec0_10_io_parallelOutput_9,{bufferVec0_10_io_parallelOutput_8,{bufferVec0_10_io_parallelOutput_7,{bufferVec0_10_io_parallelOutput_6,{bufferVec0_10_io_parallelOutput_5,{bufferVec0_10_io_parallelOutput_4,{bufferVec0_10_io_parallelOutput_3,{bufferVec0_10_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_18,_zz__zz_io_parallelInput_0_18_1}}}}}}}}}}};
  assign bufferVec0_9_io_parallelInput_0 = _zz_io_parallelInput_0_18[254 : 0];
  assign bufferVec0_9_io_parallelInput_1 = _zz_io_parallelInput_0_18[509 : 255];
  assign bufferVec0_9_io_parallelInput_2 = _zz_io_parallelInput_0_18[764 : 510];
  assign bufferVec0_9_io_parallelInput_3 = _zz_io_parallelInput_0_18[1019 : 765];
  assign bufferVec0_9_io_parallelInput_4 = _zz_io_parallelInput_0_18[1274 : 1020];
  assign bufferVec0_9_io_parallelInput_5 = _zz_io_parallelInput_0_18[1529 : 1275];
  assign bufferVec0_9_io_parallelInput_6 = _zz_io_parallelInput_0_18[1784 : 1530];
  assign bufferVec0_9_io_parallelInput_7 = _zz_io_parallelInput_0_18[2039 : 1785];
  assign bufferVec0_9_io_parallelInput_8 = _zz_io_parallelInput_0_18[2294 : 2040];
  assign bufferVec0_9_io_parallelInput_9 = _zz_io_parallelInput_0_18[2549 : 2295];
  assign bufferVec0_9_io_parallelInput_10 = _zz_io_parallelInput_0_18[2804 : 2550];
  assign bufferVec0_9_io_parallelInput_11 = _zz_io_parallelInput_0_18[3059 : 2805];
  assign _zz_io_parallelInput_0_19 = {bufferVec1_10_io_parallelOutput_11,{bufferVec1_10_io_parallelOutput_10,{bufferVec1_10_io_parallelOutput_9,{bufferVec1_10_io_parallelOutput_8,{bufferVec1_10_io_parallelOutput_7,{bufferVec1_10_io_parallelOutput_6,{bufferVec1_10_io_parallelOutput_5,{bufferVec1_10_io_parallelOutput_4,{bufferVec1_10_io_parallelOutput_3,{bufferVec1_10_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_19,_zz__zz_io_parallelInput_0_19_1}}}}}}}}}}};
  assign bufferVec1_9_io_parallelInput_0 = _zz_io_parallelInput_0_19[254 : 0];
  assign bufferVec1_9_io_parallelInput_1 = _zz_io_parallelInput_0_19[509 : 255];
  assign bufferVec1_9_io_parallelInput_2 = _zz_io_parallelInput_0_19[764 : 510];
  assign bufferVec1_9_io_parallelInput_3 = _zz_io_parallelInput_0_19[1019 : 765];
  assign bufferVec1_9_io_parallelInput_4 = _zz_io_parallelInput_0_19[1274 : 1020];
  assign bufferVec1_9_io_parallelInput_5 = _zz_io_parallelInput_0_19[1529 : 1275];
  assign bufferVec1_9_io_parallelInput_6 = _zz_io_parallelInput_0_19[1784 : 1530];
  assign bufferVec1_9_io_parallelInput_7 = _zz_io_parallelInput_0_19[2039 : 1785];
  assign bufferVec1_9_io_parallelInput_8 = _zz_io_parallelInput_0_19[2294 : 2040];
  assign bufferVec1_9_io_parallelInput_9 = _zz_io_parallelInput_0_19[2549 : 2295];
  assign bufferVec1_9_io_parallelInput_10 = _zz_io_parallelInput_0_19[2804 : 2550];
  assign bufferVec1_9_io_parallelInput_11 = _zz_io_parallelInput_0_19[3059 : 2805];
  assign _zz_io_parallelInput_0_20 = {bufferVec0_11_io_parallelOutput_11,{bufferVec0_11_io_parallelOutput_10,{bufferVec0_11_io_parallelOutput_9,{bufferVec0_11_io_parallelOutput_8,{bufferVec0_11_io_parallelOutput_7,{bufferVec0_11_io_parallelOutput_6,{bufferVec0_11_io_parallelOutput_5,{bufferVec0_11_io_parallelOutput_4,{bufferVec0_11_io_parallelOutput_3,{bufferVec0_11_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_20,_zz__zz_io_parallelInput_0_20_1}}}}}}}}}}};
  assign bufferVec0_10_io_parallelInput_0 = _zz_io_parallelInput_0_20[254 : 0];
  assign bufferVec0_10_io_parallelInput_1 = _zz_io_parallelInput_0_20[509 : 255];
  assign bufferVec0_10_io_parallelInput_2 = _zz_io_parallelInput_0_20[764 : 510];
  assign bufferVec0_10_io_parallelInput_3 = _zz_io_parallelInput_0_20[1019 : 765];
  assign bufferVec0_10_io_parallelInput_4 = _zz_io_parallelInput_0_20[1274 : 1020];
  assign bufferVec0_10_io_parallelInput_5 = _zz_io_parallelInput_0_20[1529 : 1275];
  assign bufferVec0_10_io_parallelInput_6 = _zz_io_parallelInput_0_20[1784 : 1530];
  assign bufferVec0_10_io_parallelInput_7 = _zz_io_parallelInput_0_20[2039 : 1785];
  assign bufferVec0_10_io_parallelInput_8 = _zz_io_parallelInput_0_20[2294 : 2040];
  assign bufferVec0_10_io_parallelInput_9 = _zz_io_parallelInput_0_20[2549 : 2295];
  assign bufferVec0_10_io_parallelInput_10 = _zz_io_parallelInput_0_20[2804 : 2550];
  assign bufferVec0_10_io_parallelInput_11 = _zz_io_parallelInput_0_20[3059 : 2805];
  assign _zz_io_parallelInput_0_21 = {bufferVec1_11_io_parallelOutput_11,{bufferVec1_11_io_parallelOutput_10,{bufferVec1_11_io_parallelOutput_9,{bufferVec1_11_io_parallelOutput_8,{bufferVec1_11_io_parallelOutput_7,{bufferVec1_11_io_parallelOutput_6,{bufferVec1_11_io_parallelOutput_5,{bufferVec1_11_io_parallelOutput_4,{bufferVec1_11_io_parallelOutput_3,{bufferVec1_11_io_parallelOutput_2,{_zz__zz_io_parallelInput_0_21,_zz__zz_io_parallelInput_0_21_1}}}}}}}}}}};
  assign bufferVec1_10_io_parallelInput_0 = _zz_io_parallelInput_0_21[254 : 0];
  assign bufferVec1_10_io_parallelInput_1 = _zz_io_parallelInput_0_21[509 : 255];
  assign bufferVec1_10_io_parallelInput_2 = _zz_io_parallelInput_0_21[764 : 510];
  assign bufferVec1_10_io_parallelInput_3 = _zz_io_parallelInput_0_21[1019 : 765];
  assign bufferVec1_10_io_parallelInput_4 = _zz_io_parallelInput_0_21[1274 : 1020];
  assign bufferVec1_10_io_parallelInput_5 = _zz_io_parallelInput_0_21[1529 : 1275];
  assign bufferVec1_10_io_parallelInput_6 = _zz_io_parallelInput_0_21[1784 : 1530];
  assign bufferVec1_10_io_parallelInput_7 = _zz_io_parallelInput_0_21[2039 : 1785];
  assign bufferVec1_10_io_parallelInput_8 = _zz_io_parallelInput_0_21[2294 : 2040];
  assign bufferVec1_10_io_parallelInput_9 = _zz_io_parallelInput_0_21[2549 : 2295];
  assign bufferVec1_10_io_parallelInput_10 = _zz_io_parallelInput_0_21[2804 : 2550];
  assign bufferVec1_10_io_parallelInput_11 = _zz_io_parallelInput_0_21[3059 : 2805];
  assign _zz_io_parallelInput_0_22 = 3060'h0;
  assign bufferVec0_11_io_parallelInput_0 = _zz_io_parallelInput_0_22[254 : 0];
  assign bufferVec0_11_io_parallelInput_1 = _zz_io_parallelInput_0_22[509 : 255];
  assign bufferVec0_11_io_parallelInput_2 = _zz_io_parallelInput_0_22[764 : 510];
  assign bufferVec0_11_io_parallelInput_3 = _zz_io_parallelInput_0_22[1019 : 765];
  assign bufferVec0_11_io_parallelInput_4 = _zz_io_parallelInput_0_22[1274 : 1020];
  assign bufferVec0_11_io_parallelInput_5 = _zz_io_parallelInput_0_22[1529 : 1275];
  assign bufferVec0_11_io_parallelInput_6 = _zz_io_parallelInput_0_22[1784 : 1530];
  assign bufferVec0_11_io_parallelInput_7 = _zz_io_parallelInput_0_22[2039 : 1785];
  assign bufferVec0_11_io_parallelInput_8 = _zz_io_parallelInput_0_22[2294 : 2040];
  assign bufferVec0_11_io_parallelInput_9 = _zz_io_parallelInput_0_22[2549 : 2295];
  assign bufferVec0_11_io_parallelInput_10 = _zz_io_parallelInput_0_22[2804 : 2550];
  assign bufferVec0_11_io_parallelInput_11 = _zz_io_parallelInput_0_22[3059 : 2805];
  assign _zz_io_parallelInput_0_23 = 3060'h0;
  assign bufferVec1_11_io_parallelInput_0 = _zz_io_parallelInput_0_23[254 : 0];
  assign bufferVec1_11_io_parallelInput_1 = _zz_io_parallelInput_0_23[509 : 255];
  assign bufferVec1_11_io_parallelInput_2 = _zz_io_parallelInput_0_23[764 : 510];
  assign bufferVec1_11_io_parallelInput_3 = _zz_io_parallelInput_0_23[1019 : 765];
  assign bufferVec1_11_io_parallelInput_4 = _zz_io_parallelInput_0_23[1274 : 1020];
  assign bufferVec1_11_io_parallelInput_5 = _zz_io_parallelInput_0_23[1529 : 1275];
  assign bufferVec1_11_io_parallelInput_6 = _zz_io_parallelInput_0_23[1784 : 1530];
  assign bufferVec1_11_io_parallelInput_7 = _zz_io_parallelInput_0_23[2039 : 1785];
  assign bufferVec1_11_io_parallelInput_8 = _zz_io_parallelInput_0_23[2294 : 2040];
  assign bufferVec1_11_io_parallelInput_9 = _zz_io_parallelInput_0_23[2549 : 2295];
  assign bufferVec1_11_io_parallelInput_10 = _zz_io_parallelInput_0_23[2804 : 2550];
  assign bufferVec1_11_io_parallelInput_11 = _zz_io_parallelInput_0_23[3059 : 2805];
  assign fsm_wantExit = 1'b0;
  always @(*) begin
    fsm_wantStart = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
      end
      fsm_enumDef_1_R0T1 : begin
      end
      default : begin
        fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign fsm_wantKill = 1'b0;
  always @(*) begin
    io_output_valid = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_valid = 1'b1;
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_valid = 1'b1;
      end
      default : begin
      end
    endcase
  end

  assign _zz_io_output_payload_stateElements_0 = 3060'h0;
  always @(*) begin
    io_output_payload_stateElements_0 = _zz_io_output_payload_stateElements_0[254 : 0];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_0 = _zz_io_output_payload_stateElements_0_1[254 : 0];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_0 = _zz_io_output_payload_stateElements_0_2[254 : 0];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_1 = _zz_io_output_payload_stateElements_0[509 : 255];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_1 = _zz_io_output_payload_stateElements_0_1[509 : 255];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_1 = _zz_io_output_payload_stateElements_0_2[509 : 255];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_2 = _zz_io_output_payload_stateElements_0[764 : 510];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_2 = _zz_io_output_payload_stateElements_0_1[764 : 510];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_2 = _zz_io_output_payload_stateElements_0_2[764 : 510];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_3 = _zz_io_output_payload_stateElements_0[1019 : 765];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_3 = _zz_io_output_payload_stateElements_0_1[1019 : 765];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_3 = _zz_io_output_payload_stateElements_0_2[1019 : 765];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_4 = _zz_io_output_payload_stateElements_0[1274 : 1020];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_4 = _zz_io_output_payload_stateElements_0_1[1274 : 1020];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_4 = _zz_io_output_payload_stateElements_0_2[1274 : 1020];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_5 = _zz_io_output_payload_stateElements_0[1529 : 1275];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_5 = _zz_io_output_payload_stateElements_0_1[1529 : 1275];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_5 = _zz_io_output_payload_stateElements_0_2[1529 : 1275];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_6 = _zz_io_output_payload_stateElements_0[1784 : 1530];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_6 = _zz_io_output_payload_stateElements_0_1[1784 : 1530];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_6 = _zz_io_output_payload_stateElements_0_2[1784 : 1530];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_7 = _zz_io_output_payload_stateElements_0[2039 : 1785];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_7 = _zz_io_output_payload_stateElements_0_1[2039 : 1785];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_7 = _zz_io_output_payload_stateElements_0_2[2039 : 1785];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_8 = _zz_io_output_payload_stateElements_0[2294 : 2040];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_8 = _zz_io_output_payload_stateElements_0_1[2294 : 2040];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_8 = _zz_io_output_payload_stateElements_0_2[2294 : 2040];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_9 = _zz_io_output_payload_stateElements_0[2549 : 2295];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_9 = _zz_io_output_payload_stateElements_0_1[2549 : 2295];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_9 = _zz_io_output_payload_stateElements_0_2[2549 : 2295];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_10 = _zz_io_output_payload_stateElements_0[2804 : 2550];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_10 = _zz_io_output_payload_stateElements_0_1[2804 : 2550];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_10 = _zz_io_output_payload_stateElements_0_2[2804 : 2550];
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    io_output_payload_stateElements_11 = _zz_io_output_payload_stateElements_0[3059 : 2805];
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        io_output_payload_stateElements_11 = _zz_io_output_payload_stateElements_0_1[3059 : 2805];
      end
      fsm_enumDef_1_R0T1 : begin
        io_output_payload_stateElements_11 = _zz_io_output_payload_stateElements_0_2[3059 : 2805];
      end
      default : begin
      end
    endcase
  end

  assign io_output_payload_isFull = fsm_outContext_isFull;
  assign io_output_payload_fullRound = fsm_outContext_fullRound;
  assign io_output_payload_partialRound = fsm_outContext_partialRound;
  assign io_output_payload_stateSize = fsm_outContext_stateSize;
  assign io_output_payload_stateID = fsm_outContext_stateID;
  always @(*) begin
    bufferEna0 = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
        if(io_input_valid) begin
          bufferEna0 = 1'b1;
        end
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
      end
      fsm_enumDef_1_R0T1 : begin
        if(io_input_valid) begin
          bufferEna0 = 1'b1;
        end
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bufferEna1 = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
        if(io_input_valid) begin
          bufferEna1 = 1'b1;
        end
      end
      fsm_enumDef_1_T0R1 : begin
        if(io_input_valid) begin
          bufferEna1 = 1'b1;
        end
      end
      fsm_enumDef_1_R0T1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bufferInit0 = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
        bufferInit0 = 1'b1;
      end
      fsm_enumDef_1_R0T1 : begin
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    bufferInit1 = 1'b0;
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
      end
      fsm_enumDef_1_R1R0 : begin
      end
      fsm_enumDef_1_T0R1 : begin
      end
      fsm_enumDef_1_R0T1 : begin
        bufferInit1 = 1'b1;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    fsm_stateNext = fsm_stateReg;
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
        if(io_input_valid) begin
          if(when_MDSMatrixAdders_l257) begin
            fsm_stateNext = fsm_enumDef_1_T0R1;
          end
        end
      end
      fsm_enumDef_1_R1R0 : begin
        if(io_input_valid) begin
          if(when_MDSMatrixAdders_l270) begin
            fsm_stateNext = fsm_enumDef_1_R0T1;
          end
        end
      end
      fsm_enumDef_1_T0R1 : begin
        if(when_MDSMatrixAdders_l292) begin
          fsm_stateNext = fsm_enumDef_1_R0T1;
        end else begin
          if(when_MDSMatrixAdders_l296) begin
            fsm_stateNext = fsm_enumDef_1_R1R0;
          end
        end
      end
      fsm_enumDef_1_R0T1 : begin
        if(when_MDSMatrixAdders_l317) begin
          fsm_stateNext = fsm_enumDef_1_T0R1;
        end else begin
          if(when_MDSMatrixAdders_l321) begin
            fsm_stateNext = fsm_enumDef_1_R0R1;
          end
        end
      end
      default : begin
      end
    endcase
    if(fsm_wantStart) begin
      fsm_stateNext = fsm_enumDef_1_R0R1;
    end
    if(fsm_wantKill) begin
      fsm_stateNext = fsm_enumDef_1_BOOT;
    end
  end

  assign when_MDSMatrixAdders_l257 = (fsm_inCount == _zz_when_MDSMatrixAdders_l257);
  assign when_MDSMatrixAdders_l270 = (fsm_inCount == _zz_when_MDSMatrixAdders_l270);
  assign _zz_io_output_payload_stateElements_0_1 = {bufferVec0_0_io_parallelOutput_11,{bufferVec0_0_io_parallelOutput_10,{bufferVec0_0_io_parallelOutput_9,{bufferVec0_0_io_parallelOutput_8,{bufferVec0_0_io_parallelOutput_7,{bufferVec0_0_io_parallelOutput_6,{bufferVec0_0_io_parallelOutput_5,{bufferVec0_0_io_parallelOutput_4,{bufferVec0_0_io_parallelOutput_3,{bufferVec0_0_io_parallelOutput_2,{_zz__zz_io_output_payload_stateElements_0_1,_zz__zz_io_output_payload_stateElements_0_1_1}}}}}}}}}}};
  assign when_MDSMatrixAdders_l292 = (io_input_valid && (fsm_inCount == _zz_when_MDSMatrixAdders_l292));
  assign when_MDSMatrixAdders_l296 = (fsm_outCount == _zz_when_MDSMatrixAdders_l296);
  assign _zz_io_output_payload_stateElements_0_2 = {bufferVec1_0_io_parallelOutput_11,{bufferVec1_0_io_parallelOutput_10,{bufferVec1_0_io_parallelOutput_9,{bufferVec1_0_io_parallelOutput_8,{bufferVec1_0_io_parallelOutput_7,{bufferVec1_0_io_parallelOutput_6,{bufferVec1_0_io_parallelOutput_5,{bufferVec1_0_io_parallelOutput_4,{bufferVec1_0_io_parallelOutput_3,{bufferVec1_0_io_parallelOutput_2,{_zz__zz_io_output_payload_stateElements_0_2,_zz__zz_io_output_payload_stateElements_0_2_1}}}}}}}}}}};
  assign when_MDSMatrixAdders_l317 = (io_input_valid && (fsm_inCount == _zz_when_MDSMatrixAdders_l317));
  assign when_MDSMatrixAdders_l321 = (fsm_outCount == _zz_when_MDSMatrixAdders_l321);
  assign when_StateMachine_l222 = ((fsm_stateReg == fsm_enumDef_1_R0R1) && (! (fsm_stateNext == fsm_enumDef_1_R0R1)));
  assign when_StateMachine_l222_1 = ((fsm_stateReg == fsm_enumDef_1_R1R0) && (! (fsm_stateNext == fsm_enumDef_1_R1R0)));
  assign when_StateMachine_l222_2 = ((fsm_stateReg == fsm_enumDef_1_T0R1) && (! (fsm_stateNext == fsm_enumDef_1_T0R1)));
  assign when_StateMachine_l222_3 = ((fsm_stateReg == fsm_enumDef_1_R0T1) && (! (fsm_stateNext == fsm_enumDef_1_R0T1)));
  always @(posedge clk) begin
    if(!resetn) begin
      fsm_inCount <= 4'b0000;
      fsm_outCount <= 4'b0000;
      fsm_stateReg <= fsm_enumDef_1_BOOT;
    end else begin
      fsm_stateReg <= fsm_stateNext;
      case(fsm_stateReg)
        fsm_enumDef_1_R0R1 : begin
          if(io_input_valid) begin
            fsm_inCount <= (fsm_inCount + 4'b0001);
          end
        end
        fsm_enumDef_1_R1R0 : begin
          if(io_input_valid) begin
            fsm_inCount <= (fsm_inCount + 4'b0001);
          end
        end
        fsm_enumDef_1_T0R1 : begin
          fsm_outCount <= (fsm_outCount + 4'b0001);
          if(io_input_valid) begin
            fsm_inCount <= (fsm_inCount + 4'b0001);
          end
          if(when_MDSMatrixAdders_l292) begin
            fsm_inCount <= 4'b0000;
          end
        end
        fsm_enumDef_1_R0T1 : begin
          fsm_outCount <= (fsm_outCount + 4'b0001);
          if(io_input_valid) begin
            fsm_inCount <= (fsm_inCount + 4'b0001);
          end
          if(when_MDSMatrixAdders_l317) begin
            fsm_inCount <= 4'b0000;
          end
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l222) begin
        fsm_inCount <= 4'b0000;
      end
      if(when_StateMachine_l222_1) begin
        fsm_inCount <= 4'b0000;
      end
      if(when_StateMachine_l222_2) begin
        fsm_outCount <= 4'b0000;
      end
      if(when_StateMachine_l222_3) begin
        fsm_outCount <= 4'b0000;
      end
    end
  end

  always @(posedge clk) begin
    case(fsm_stateReg)
      fsm_enumDef_1_R0R1 : begin
        if(io_input_valid) begin
          if(when_MDSMatrixAdders_l257) begin
            fsm_outContext_isFull <= io_input_payload_isFull;
            fsm_outContext_fullRound <= io_input_payload_fullRound;
            fsm_outContext_partialRound <= io_input_payload_partialRound;
            fsm_outContext_stateSize <= io_input_payload_stateSize;
            fsm_outContext_stateID <= io_input_payload_stateID;
          end
        end
      end
      fsm_enumDef_1_R1R0 : begin
        if(io_input_valid) begin
          if(when_MDSMatrixAdders_l270) begin
            fsm_outContext_isFull <= io_input_payload_isFull;
            fsm_outContext_fullRound <= io_input_payload_fullRound;
            fsm_outContext_partialRound <= io_input_payload_partialRound;
            fsm_outContext_stateSize <= io_input_payload_stateSize;
            fsm_outContext_stateID <= io_input_payload_stateID;
          end
        end
      end
      fsm_enumDef_1_T0R1 : begin
        if(when_MDSMatrixAdders_l292) begin
          fsm_outContext_isFull <= io_input_payload_isFull;
          fsm_outContext_fullRound <= io_input_payload_fullRound;
          fsm_outContext_partialRound <= io_input_payload_partialRound;
          fsm_outContext_stateSize <= io_input_payload_stateSize;
          fsm_outContext_stateID <= io_input_payload_stateID;
        end
      end
      fsm_enumDef_1_R0T1 : begin
        if(when_MDSMatrixAdders_l317) begin
          fsm_outContext_isFull <= io_input_payload_isFull;
          fsm_outContext_fullRound <= io_input_payload_fullRound;
          fsm_outContext_partialRound <= io_input_payload_partialRound;
          fsm_outContext_stateSize <= io_input_payload_stateSize;
          fsm_outContext_stateID <= io_input_payload_stateID;
        end
      end
      default : begin
      end
    endcase
  end


endmodule

module AdderTree (
  input               io_input_valid,
  input      [254:0]  io_input_payload_0,
  input      [254:0]  io_input_payload_1,
  input      [254:0]  io_input_payload_2,
  input      [254:0]  io_input_payload_3,
  input      [254:0]  io_input_payload_4,
  input      [254:0]  io_input_payload_5,
  input      [254:0]  io_input_payload_6,
  input      [254:0]  io_input_payload_7,
  input      [254:0]  io_input_payload_8,
  input      [254:0]  io_input_payload_9,
  input      [254:0]  io_input_payload_10,
  input      [254:0]  io_input_payload_11,
  output              io_output_valid,
  output     [254:0]  io_output_payload,
  input               clk,
  input               resetn
);

  wire       [254:0]  modAdderPiped_28_io_op1;
  wire       [254:0]  modAdderPiped_28_io_op2;
  wire       [254:0]  modAdderPiped_29_io_op1;
  wire       [254:0]  modAdderPiped_29_io_op2;
  wire       [254:0]  modAdderPiped_30_io_op1;
  wire       [254:0]  modAdderPiped_30_io_op2;
  wire       [254:0]  modAdderPiped_31_io_op1;
  wire       [254:0]  modAdderPiped_31_io_op2;
  wire       [254:0]  modAdderPiped_32_io_op1;
  wire       [254:0]  modAdderPiped_32_io_op2;
  wire       [254:0]  modAdderPiped_22_io_res;
  wire       [254:0]  modAdderPiped_23_io_res;
  wire       [254:0]  modAdderPiped_24_io_res;
  wire       [254:0]  modAdderPiped_25_io_res;
  wire       [254:0]  modAdderPiped_26_io_res;
  wire       [254:0]  modAdderPiped_27_io_res;
  wire       [254:0]  modAdderPiped_28_io_res;
  wire       [254:0]  modAdderPiped_29_io_res;
  wire       [254:0]  modAdderPiped_30_io_res;
  wire       [254:0]  modAdderPiped_31_io_res;
  wire       [254:0]  modAdderPiped_32_io_res;
  wire       [1529:0] _zz_io_op1;
  wire       [764:0]  _zz_io_op1_1;
  reg        [254:0]  _zz_io_op1_2;
  reg        [254:0]  _zz_io_op1_3;
  reg        [254:0]  _zz_io_op1_4;
  reg        [254:0]  _zz_io_op1_5;
  reg        [254:0]  _zz_io_op1_6;
  reg        [254:0]  _zz_io_op1_7;
  reg        [254:0]  _zz_io_op1_8;
  reg        [254:0]  _zz_io_op1_9;
  reg        [254:0]  _zz_io_op1_10;
  reg        [254:0]  _zz_io_op1_11;
  reg        [254:0]  _zz_io_op1_12;
  reg        [254:0]  _zz_io_op1_13;
  reg        [254:0]  _zz_io_op1_14;
  reg        [254:0]  _zz_io_op1_15;
  reg        [254:0]  _zz_io_op1_16;
  reg        [254:0]  _zz_io_op1_17;
  wire       [509:0]  _zz_io_op1_18;
  reg                 io_input_valid_delay_1;
  reg                 io_input_valid_delay_2;
  reg                 io_input_valid_delay_3;
  reg                 io_input_valid_delay_4;
  reg                 io_input_valid_delay_5;
  reg                 io_input_valid_delay_6;
  reg                 io_input_valid_delay_7;
  reg                 io_input_valid_delay_8;
  reg                 io_input_valid_delay_9;
  reg                 io_input_valid_delay_10;
  reg                 io_input_valid_delay_11;
  reg                 io_input_valid_delay_12;
  reg                 io_input_valid_delay_13;
  reg                 io_input_valid_delay_14;
  reg                 io_input_valid_delay_15;
  reg                 io_input_valid_delay_16;
  reg                 io_input_valid_delay_17;
  reg                 io_input_valid_delay_18;
  reg                 io_input_valid_delay_19;
  reg                 io_input_valid_delay_20;
  reg                 io_input_valid_delay_21;
  reg                 io_input_valid_delay_22;
  reg                 io_input_valid_delay_23;
  reg                 io_input_valid_delay_24;
  reg                 io_input_valid_delay_25;
  reg                 io_input_valid_delay_26;
  reg                 io_input_valid_delay_27;
  reg                 io_input_valid_delay_28;
  reg                 io_input_valid_delay_29;
  reg                 io_input_valid_delay_30;
  reg                 io_input_valid_delay_31;
  reg                 io_input_valid_delay_32;
  reg                 io_input_valid_delay_33;
  reg                 io_input_valid_delay_34;
  reg                 io_input_valid_delay_35;
  reg                 io_input_valid_delay_36;
  reg                 io_input_valid_delay_37;
  reg                 io_input_valid_delay_38;
  reg                 io_input_valid_delay_39;
  reg                 io_input_valid_delay_40;
  reg                 io_input_valid_delay_41;
  reg                 io_input_valid_delay_42;
  reg                 io_input_valid_delay_43;
  reg                 io_input_valid_delay_44;
  reg                 io_input_valid_delay_45;
  reg                 io_input_valid_delay_46;
  reg                 io_input_valid_delay_47;
  reg                 io_input_valid_delay_48;
  reg                 io_input_valid_delay_49;
  reg                 io_input_valid_delay_50;
  reg                 io_input_valid_delay_51;
  reg                 io_input_valid_delay_52;
  reg                 io_input_valid_delay_53;
  reg                 io_input_valid_delay_54;
  reg                 io_input_valid_delay_55;
  reg                 io_input_valid_delay_56;
  reg                 io_input_valid_delay_57;
  reg                 io_input_valid_delay_58;
  reg                 io_input_valid_delay_59;
  reg                 io_input_valid_delay_60;
  reg                 io_input_valid_delay_61;
  reg                 io_input_valid_delay_62;
  reg                 io_input_valid_delay_63;
  reg                 io_input_valid_delay_64;

  ModAdderPiped modAdderPiped_22 (
    .io_op1    (io_input_payload_0[254:0]       ), //i
    .io_op2    (io_input_payload_1[254:0]       ), //i
    .io_res    (modAdderPiped_22_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_23 (
    .io_op1    (io_input_payload_2[254:0]       ), //i
    .io_op2    (io_input_payload_3[254:0]       ), //i
    .io_res    (modAdderPiped_23_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_24 (
    .io_op1    (io_input_payload_4[254:0]       ), //i
    .io_op2    (io_input_payload_5[254:0]       ), //i
    .io_res    (modAdderPiped_24_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_25 (
    .io_op1    (io_input_payload_6[254:0]       ), //i
    .io_op2    (io_input_payload_7[254:0]       ), //i
    .io_res    (modAdderPiped_25_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_26 (
    .io_op1    (io_input_payload_8[254:0]       ), //i
    .io_op2    (io_input_payload_9[254:0]       ), //i
    .io_res    (modAdderPiped_26_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_27 (
    .io_op1    (io_input_payload_10[254:0]      ), //i
    .io_op2    (io_input_payload_11[254:0]      ), //i
    .io_res    (modAdderPiped_27_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_28 (
    .io_op1    (modAdderPiped_28_io_op1[254:0]  ), //i
    .io_op2    (modAdderPiped_28_io_op2[254:0]  ), //i
    .io_res    (modAdderPiped_28_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_29 (
    .io_op1    (modAdderPiped_29_io_op1[254:0]  ), //i
    .io_op2    (modAdderPiped_29_io_op2[254:0]  ), //i
    .io_res    (modAdderPiped_29_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_30 (
    .io_op1    (modAdderPiped_30_io_op1[254:0]  ), //i
    .io_op2    (modAdderPiped_30_io_op2[254:0]  ), //i
    .io_res    (modAdderPiped_30_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_31 (
    .io_op1    (modAdderPiped_31_io_op1[254:0]  ), //i
    .io_op2    (modAdderPiped_31_io_op2[254:0]  ), //i
    .io_res    (modAdderPiped_31_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  ModAdderPiped modAdderPiped_32 (
    .io_op1    (modAdderPiped_32_io_op1[254:0]  ), //i
    .io_op2    (modAdderPiped_32_io_op2[254:0]  ), //i
    .io_res    (modAdderPiped_32_io_res[254:0]  ), //o
    .clk       (clk                             ), //i
    .resetn    (resetn                          )  //i
  );
  assign _zz_io_op1 = {modAdderPiped_27_io_res,{modAdderPiped_26_io_res,{modAdderPiped_25_io_res,{modAdderPiped_24_io_res,{modAdderPiped_23_io_res,modAdderPiped_22_io_res}}}}};
  assign modAdderPiped_28_io_op1 = _zz_io_op1[254 : 0];
  assign modAdderPiped_28_io_op2 = _zz_io_op1[509 : 255];
  assign modAdderPiped_29_io_op1 = _zz_io_op1[764 : 510];
  assign modAdderPiped_29_io_op2 = _zz_io_op1[1019 : 765];
  assign modAdderPiped_30_io_op1 = _zz_io_op1[1274 : 1020];
  assign modAdderPiped_30_io_op2 = _zz_io_op1[1529 : 1275];
  assign _zz_io_op1_1 = {modAdderPiped_30_io_res,{modAdderPiped_29_io_res,modAdderPiped_28_io_res}};
  assign modAdderPiped_31_io_op1 = _zz_io_op1_1[254 : 0];
  assign modAdderPiped_31_io_op2 = _zz_io_op1_1[509 : 255];
  assign _zz_io_op1_18 = {_zz_io_op1_17,modAdderPiped_31_io_res};
  assign modAdderPiped_32_io_op1 = _zz_io_op1_18[254 : 0];
  assign modAdderPiped_32_io_op2 = _zz_io_op1_18[509 : 255];
  assign io_output_valid = io_input_valid_delay_64;
  assign io_output_payload = modAdderPiped_32_io_res;
  always @(posedge clk) begin
    _zz_io_op1_2 <= _zz_io_op1_1[764 : 510];
    _zz_io_op1_3 <= _zz_io_op1_2;
    _zz_io_op1_4 <= _zz_io_op1_3;
    _zz_io_op1_5 <= _zz_io_op1_4;
    _zz_io_op1_6 <= _zz_io_op1_5;
    _zz_io_op1_7 <= _zz_io_op1_6;
    _zz_io_op1_8 <= _zz_io_op1_7;
    _zz_io_op1_9 <= _zz_io_op1_8;
    _zz_io_op1_10 <= _zz_io_op1_9;
    _zz_io_op1_11 <= _zz_io_op1_10;
    _zz_io_op1_12 <= _zz_io_op1_11;
    _zz_io_op1_13 <= _zz_io_op1_12;
    _zz_io_op1_14 <= _zz_io_op1_13;
    _zz_io_op1_15 <= _zz_io_op1_14;
    _zz_io_op1_16 <= _zz_io_op1_15;
    _zz_io_op1_17 <= _zz_io_op1_16;
  end

  always @(posedge clk) begin
    if(!resetn) begin
      io_input_valid_delay_1 <= 1'b0;
      io_input_valid_delay_2 <= 1'b0;
      io_input_valid_delay_3 <= 1'b0;
      io_input_valid_delay_4 <= 1'b0;
      io_input_valid_delay_5 <= 1'b0;
      io_input_valid_delay_6 <= 1'b0;
      io_input_valid_delay_7 <= 1'b0;
      io_input_valid_delay_8 <= 1'b0;
      io_input_valid_delay_9 <= 1'b0;
      io_input_valid_delay_10 <= 1'b0;
      io_input_valid_delay_11 <= 1'b0;
      io_input_valid_delay_12 <= 1'b0;
      io_input_valid_delay_13 <= 1'b0;
      io_input_valid_delay_14 <= 1'b0;
      io_input_valid_delay_15 <= 1'b0;
      io_input_valid_delay_16 <= 1'b0;
      io_input_valid_delay_17 <= 1'b0;
      io_input_valid_delay_18 <= 1'b0;
      io_input_valid_delay_19 <= 1'b0;
      io_input_valid_delay_20 <= 1'b0;
      io_input_valid_delay_21 <= 1'b0;
      io_input_valid_delay_22 <= 1'b0;
      io_input_valid_delay_23 <= 1'b0;
      io_input_valid_delay_24 <= 1'b0;
      io_input_valid_delay_25 <= 1'b0;
      io_input_valid_delay_26 <= 1'b0;
      io_input_valid_delay_27 <= 1'b0;
      io_input_valid_delay_28 <= 1'b0;
      io_input_valid_delay_29 <= 1'b0;
      io_input_valid_delay_30 <= 1'b0;
      io_input_valid_delay_31 <= 1'b0;
      io_input_valid_delay_32 <= 1'b0;
      io_input_valid_delay_33 <= 1'b0;
      io_input_valid_delay_34 <= 1'b0;
      io_input_valid_delay_35 <= 1'b0;
      io_input_valid_delay_36 <= 1'b0;
      io_input_valid_delay_37 <= 1'b0;
      io_input_valid_delay_38 <= 1'b0;
      io_input_valid_delay_39 <= 1'b0;
      io_input_valid_delay_40 <= 1'b0;
      io_input_valid_delay_41 <= 1'b0;
      io_input_valid_delay_42 <= 1'b0;
      io_input_valid_delay_43 <= 1'b0;
      io_input_valid_delay_44 <= 1'b0;
      io_input_valid_delay_45 <= 1'b0;
      io_input_valid_delay_46 <= 1'b0;
      io_input_valid_delay_47 <= 1'b0;
      io_input_valid_delay_48 <= 1'b0;
      io_input_valid_delay_49 <= 1'b0;
      io_input_valid_delay_50 <= 1'b0;
      io_input_valid_delay_51 <= 1'b0;
      io_input_valid_delay_52 <= 1'b0;
      io_input_valid_delay_53 <= 1'b0;
      io_input_valid_delay_54 <= 1'b0;
      io_input_valid_delay_55 <= 1'b0;
      io_input_valid_delay_56 <= 1'b0;
      io_input_valid_delay_57 <= 1'b0;
      io_input_valid_delay_58 <= 1'b0;
      io_input_valid_delay_59 <= 1'b0;
      io_input_valid_delay_60 <= 1'b0;
      io_input_valid_delay_61 <= 1'b0;
      io_input_valid_delay_62 <= 1'b0;
      io_input_valid_delay_63 <= 1'b0;
      io_input_valid_delay_64 <= 1'b0;
    end else begin
      io_input_valid_delay_1 <= io_input_valid;
      io_input_valid_delay_2 <= io_input_valid_delay_1;
      io_input_valid_delay_3 <= io_input_valid_delay_2;
      io_input_valid_delay_4 <= io_input_valid_delay_3;
      io_input_valid_delay_5 <= io_input_valid_delay_4;
      io_input_valid_delay_6 <= io_input_valid_delay_5;
      io_input_valid_delay_7 <= io_input_valid_delay_6;
      io_input_valid_delay_8 <= io_input_valid_delay_7;
      io_input_valid_delay_9 <= io_input_valid_delay_8;
      io_input_valid_delay_10 <= io_input_valid_delay_9;
      io_input_valid_delay_11 <= io_input_valid_delay_10;
      io_input_valid_delay_12 <= io_input_valid_delay_11;
      io_input_valid_delay_13 <= io_input_valid_delay_12;
      io_input_valid_delay_14 <= io_input_valid_delay_13;
      io_input_valid_delay_15 <= io_input_valid_delay_14;
      io_input_valid_delay_16 <= io_input_valid_delay_15;
      io_input_valid_delay_17 <= io_input_valid_delay_16;
      io_input_valid_delay_18 <= io_input_valid_delay_17;
      io_input_valid_delay_19 <= io_input_valid_delay_18;
      io_input_valid_delay_20 <= io_input_valid_delay_19;
      io_input_valid_delay_21 <= io_input_valid_delay_20;
      io_input_valid_delay_22 <= io_input_valid_delay_21;
      io_input_valid_delay_23 <= io_input_valid_delay_22;
      io_input_valid_delay_24 <= io_input_valid_delay_23;
      io_input_valid_delay_25 <= io_input_valid_delay_24;
      io_input_valid_delay_26 <= io_input_valid_delay_25;
      io_input_valid_delay_27 <= io_input_valid_delay_26;
      io_input_valid_delay_28 <= io_input_valid_delay_27;
      io_input_valid_delay_29 <= io_input_valid_delay_28;
      io_input_valid_delay_30 <= io_input_valid_delay_29;
      io_input_valid_delay_31 <= io_input_valid_delay_30;
      io_input_valid_delay_32 <= io_input_valid_delay_31;
      io_input_valid_delay_33 <= io_input_valid_delay_32;
      io_input_valid_delay_34 <= io_input_valid_delay_33;
      io_input_valid_delay_35 <= io_input_valid_delay_34;
      io_input_valid_delay_36 <= io_input_valid_delay_35;
      io_input_valid_delay_37 <= io_input_valid_delay_36;
      io_input_valid_delay_38 <= io_input_valid_delay_37;
      io_input_valid_delay_39 <= io_input_valid_delay_38;
      io_input_valid_delay_40 <= io_input_valid_delay_39;
      io_input_valid_delay_41 <= io_input_valid_delay_40;
      io_input_valid_delay_42 <= io_input_valid_delay_41;
      io_input_valid_delay_43 <= io_input_valid_delay_42;
      io_input_valid_delay_44 <= io_input_valid_delay_43;
      io_input_valid_delay_45 <= io_input_valid_delay_44;
      io_input_valid_delay_46 <= io_input_valid_delay_45;
      io_input_valid_delay_47 <= io_input_valid_delay_46;
      io_input_valid_delay_48 <= io_input_valid_delay_47;
      io_input_valid_delay_49 <= io_input_valid_delay_48;
      io_input_valid_delay_50 <= io_input_valid_delay_49;
      io_input_valid_delay_51 <= io_input_valid_delay_50;
      io_input_valid_delay_52 <= io_input_valid_delay_51;
      io_input_valid_delay_53 <= io_input_valid_delay_52;
      io_input_valid_delay_54 <= io_input_valid_delay_53;
      io_input_valid_delay_55 <= io_input_valid_delay_54;
      io_input_valid_delay_56 <= io_input_valid_delay_55;
      io_input_valid_delay_57 <= io_input_valid_delay_56;
      io_input_valid_delay_58 <= io_input_valid_delay_57;
      io_input_valid_delay_59 <= io_input_valid_delay_58;
      io_input_valid_delay_60 <= io_input_valid_delay_59;
      io_input_valid_delay_61 <= io_input_valid_delay_60;
      io_input_valid_delay_62 <= io_input_valid_delay_61;
      io_input_valid_delay_63 <= io_input_valid_delay_62;
      io_input_valid_delay_64 <= io_input_valid_delay_63;
    end
  end


endmodule

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

//MontgomeryMultFlow replaced by MontgomeryMultFlow

module MontgomeryMultFlow (
  input               io_input_valid,
  input      [254:0]  io_input_payload_op1,
  input      [254:0]  io_input_payload_op2,
  output              io_output_valid,
  output     [254:0]  io_output_payload_res,
  input               clk,
  input               resetn
);

  wire                multiplierFlow_45_io_output_valid;
  wire       [509:0]  multiplierFlow_45_io_output_payload_res;
  wire                multiplierFlow_46_io_output_valid;
  wire       [511:0]  multiplierFlow_46_io_output_payload_res;
  wire                multiplierFlow_47_io_output_valid;
  wire       [511:0]  multiplierFlow_47_io_output_payload_res;
  wire       [256:0]  _zz_halfAddRes_carry;
  wire       [255:0]  _zz_adderOutput_payload_res;
  wire       [255:0]  _zz_adderOutput_payload_res_1;
  wire       [255:0]  _zz_adderOutput_payload_res_2;
  wire       [0:0]    _zz_adderOutput_payload_res_3;
  wire       [255:0]  _zz__zz_io_output_payload_res;
  wire                mulInput1_valid;
  wire       [255:0]  mulInput1_payload_op1;
  wire       [255:0]  mulInput1_payload_op2;
  wire                mulInput2_valid;
  wire       [255:0]  mulInput2_payload_op1;
  wire       [255:0]  mulInput2_payload_op2;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_1;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_2;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_3;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_4;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_5;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_6;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_7;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_8;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_9;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_10;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_11;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_12;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_13;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_14;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_15;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_16;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_17;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_18;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_19;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_20;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_21;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_22;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_23;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_24;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_25;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_26;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_27;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_28;
  reg        [509:0]  multiplierFlow_45_io_output_payload_res_delay_29;
  reg        [509:0]  mulRes0Delayed;
  wire                halfAddRes_carry;
  wire       [255:0]  halfAddRes_op1;
  wire       [253:0]  halfAddRes_op2;
  reg                 halfAdderOutput_valid;
  reg                 halfAdderOutput_payload_carry;
  reg        [255:0]  halfAdderOutput_payload_op1;
  reg        [253:0]  halfAdderOutput_payload_op2;
  reg                 adderOutput_valid;
  reg        [255:0]  adderOutput_payload_res;
  reg                 tempOutput_valid;
  reg        [255:0]  tempOutput_payload_op1;
  reg        [255:0]  tempOutput_payload_op2;
  reg                 _zz_io_output_valid;
  reg        [254:0]  _zz_io_output_payload_res;

  assign _zz_halfAddRes_carry = ({1'b0,multiplierFlow_47_io_output_payload_res[255 : 0]} + {1'b0,mulRes0Delayed[255 : 0]});
  assign _zz_adderOutput_payload_res = (halfAdderOutput_payload_op1 + _zz_adderOutput_payload_res_1);
  assign _zz_adderOutput_payload_res_1 = {2'd0, halfAdderOutput_payload_op2};
  assign _zz_adderOutput_payload_res_3 = halfAdderOutput_payload_carry;
  assign _zz_adderOutput_payload_res_2 = {255'd0, _zz_adderOutput_payload_res_3};
  assign _zz__zz_io_output_payload_res = ((tempOutput_payload_op1[255] || tempOutput_payload_op2[255]) ? tempOutput_payload_op2 : tempOutput_payload_op1);
  MultiplierFlow multiplierFlow_45 (
    .io_input_valid           (io_input_valid                                  ), //i
    .io_input_payload_op1     (io_input_payload_op1[254:0]                     ), //i
    .io_input_payload_op2     (io_input_payload_op2[254:0]                     ), //i
    .io_output_valid          (multiplierFlow_45_io_output_valid               ), //o
    .io_output_payload_res    (multiplierFlow_45_io_output_payload_res[509:0]  ), //o
    .clk                      (clk                                             ), //i
    .resetn                   (resetn                                          )  //i
  );
  MultiplierFlow_1 multiplierFlow_46 (
    .io_input_valid           (mulInput1_valid                                 ), //i
    .io_input_payload_op1     (mulInput1_payload_op1[255:0]                    ), //i
    .io_input_payload_op2     (mulInput1_payload_op2[255:0]                    ), //i
    .io_output_valid          (multiplierFlow_46_io_output_valid               ), //o
    .io_output_payload_res    (multiplierFlow_46_io_output_payload_res[511:0]  ), //o
    .clk                      (clk                                             ), //i
    .resetn                   (resetn                                          )  //i
  );
  MultiplierFlow_1 multiplierFlow_47 (
    .io_input_valid           (mulInput2_valid                                 ), //i
    .io_input_payload_op1     (mulInput2_payload_op1[255:0]                    ), //i
    .io_input_payload_op2     (mulInput2_payload_op2[255:0]                    ), //i
    .io_output_valid          (multiplierFlow_47_io_output_valid               ), //o
    .io_output_payload_res    (multiplierFlow_47_io_output_payload_res[511:0]  ), //o
    .clk                      (clk                                             ), //i
    .resetn                   (resetn                                          )  //i
  );
  assign mulInput1_valid = multiplierFlow_45_io_output_valid;
  assign mulInput1_payload_op1 = multiplierFlow_45_io_output_payload_res[255 : 0];
  assign mulInput1_payload_op2 = 256'h3d443ab0d7bf2839181b2c170004ec0653ba5bfffffe5bfdfffffffeffffffff;
  assign mulInput2_valid = multiplierFlow_46_io_output_valid;
  assign mulInput2_payload_op1 = multiplierFlow_46_io_output_payload_res[255 : 0];
  assign mulInput2_payload_op2 = 256'h73eda753299d7d483339d80809a1d80553bda402fffe5bfeffffffff00000001;
  assign halfAddRes_carry = _zz_halfAddRes_carry[256];
  assign halfAddRes_op1 = multiplierFlow_47_io_output_payload_res[511 : 256];
  assign halfAddRes_op2 = mulRes0Delayed[509 : 256];
  assign io_output_valid = _zz_io_output_valid;
  assign io_output_payload_res = _zz_io_output_payload_res;
  always @(posedge clk) begin
    multiplierFlow_45_io_output_payload_res_delay_1 <= multiplierFlow_45_io_output_payload_res;
    multiplierFlow_45_io_output_payload_res_delay_2 <= multiplierFlow_45_io_output_payload_res_delay_1;
    multiplierFlow_45_io_output_payload_res_delay_3 <= multiplierFlow_45_io_output_payload_res_delay_2;
    multiplierFlow_45_io_output_payload_res_delay_4 <= multiplierFlow_45_io_output_payload_res_delay_3;
    multiplierFlow_45_io_output_payload_res_delay_5 <= multiplierFlow_45_io_output_payload_res_delay_4;
    multiplierFlow_45_io_output_payload_res_delay_6 <= multiplierFlow_45_io_output_payload_res_delay_5;
    multiplierFlow_45_io_output_payload_res_delay_7 <= multiplierFlow_45_io_output_payload_res_delay_6;
    multiplierFlow_45_io_output_payload_res_delay_8 <= multiplierFlow_45_io_output_payload_res_delay_7;
    multiplierFlow_45_io_output_payload_res_delay_9 <= multiplierFlow_45_io_output_payload_res_delay_8;
    multiplierFlow_45_io_output_payload_res_delay_10 <= multiplierFlow_45_io_output_payload_res_delay_9;
    multiplierFlow_45_io_output_payload_res_delay_11 <= multiplierFlow_45_io_output_payload_res_delay_10;
    multiplierFlow_45_io_output_payload_res_delay_12 <= multiplierFlow_45_io_output_payload_res_delay_11;
    multiplierFlow_45_io_output_payload_res_delay_13 <= multiplierFlow_45_io_output_payload_res_delay_12;
    multiplierFlow_45_io_output_payload_res_delay_14 <= multiplierFlow_45_io_output_payload_res_delay_13;
    multiplierFlow_45_io_output_payload_res_delay_15 <= multiplierFlow_45_io_output_payload_res_delay_14;
    multiplierFlow_45_io_output_payload_res_delay_16 <= multiplierFlow_45_io_output_payload_res_delay_15;
    multiplierFlow_45_io_output_payload_res_delay_17 <= multiplierFlow_45_io_output_payload_res_delay_16;
    multiplierFlow_45_io_output_payload_res_delay_18 <= multiplierFlow_45_io_output_payload_res_delay_17;
    multiplierFlow_45_io_output_payload_res_delay_19 <= multiplierFlow_45_io_output_payload_res_delay_18;
    multiplierFlow_45_io_output_payload_res_delay_20 <= multiplierFlow_45_io_output_payload_res_delay_19;
    multiplierFlow_45_io_output_payload_res_delay_21 <= multiplierFlow_45_io_output_payload_res_delay_20;
    multiplierFlow_45_io_output_payload_res_delay_22 <= multiplierFlow_45_io_output_payload_res_delay_21;
    multiplierFlow_45_io_output_payload_res_delay_23 <= multiplierFlow_45_io_output_payload_res_delay_22;
    multiplierFlow_45_io_output_payload_res_delay_24 <= multiplierFlow_45_io_output_payload_res_delay_23;
    multiplierFlow_45_io_output_payload_res_delay_25 <= multiplierFlow_45_io_output_payload_res_delay_24;
    multiplierFlow_45_io_output_payload_res_delay_26 <= multiplierFlow_45_io_output_payload_res_delay_25;
    multiplierFlow_45_io_output_payload_res_delay_27 <= multiplierFlow_45_io_output_payload_res_delay_26;
    multiplierFlow_45_io_output_payload_res_delay_28 <= multiplierFlow_45_io_output_payload_res_delay_27;
    multiplierFlow_45_io_output_payload_res_delay_29 <= multiplierFlow_45_io_output_payload_res_delay_28;
    mulRes0Delayed <= multiplierFlow_45_io_output_payload_res_delay_29;
    halfAdderOutput_payload_carry <= halfAddRes_carry;
    halfAdderOutput_payload_op1 <= halfAddRes_op1;
    halfAdderOutput_payload_op2 <= halfAddRes_op2;
    adderOutput_payload_res <= (_zz_adderOutput_payload_res + _zz_adderOutput_payload_res_2);
    tempOutput_payload_op1 <= adderOutput_payload_res;
    tempOutput_payload_op2 <= ({1'b0,adderOutput_payload_res[254 : 0]} + {1'b0,255'h0c1258acd66282b7ccc627f7f65e27faac425bfd0001a40100000000ffffffff});
    _zz_io_output_payload_res <= _zz__zz_io_output_payload_res[254:0];
  end

  always @(posedge clk) begin
    if(!resetn) begin
      halfAdderOutput_valid <= 1'b0;
      adderOutput_valid <= 1'b0;
      tempOutput_valid <= 1'b0;
      _zz_io_output_valid <= 1'b0;
    end else begin
      halfAdderOutput_valid <= multiplierFlow_47_io_output_valid;
      adderOutput_valid <= halfAdderOutput_valid;
      tempOutput_valid <= adderOutput_valid;
      _zz_io_output_valid <= tempOutput_valid;
    end
  end


endmodule

module MDSConstantMem (
  input               io_addr_isFull,
  input      [2:0]    io_addr_fullRound,
  input      [5:0]    io_addr_partialRound,
  input      [3:0]    io_addr_stateIndex,
  input      [3:0]    io_addr_stateSize,
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  output     [254:0]  io_data_9,
  output     [254:0]  io_data_10,
  output     [254:0]  io_data_11,
  input               clk,
  input               resetn
);

  wire       [1:0]    matrixConstantMem_14_io_addr;
  wire       [2:0]    matrixConstantMem_15_io_addr;
  wire       [1:0]    matrixConstantMem_18_io_addr;
  wire       [2:0]    matrixConstantMem_19_io_addr;
  wire       [254:0]  matrixConstantMem_14_io_data_0;
  wire       [254:0]  matrixConstantMem_14_io_data_1;
  wire       [254:0]  matrixConstantMem_14_io_data_2;
  wire       [254:0]  matrixConstantMem_15_io_data_0;
  wire       [254:0]  matrixConstantMem_15_io_data_1;
  wire       [254:0]  matrixConstantMem_15_io_data_2;
  wire       [254:0]  matrixConstantMem_15_io_data_3;
  wire       [254:0]  matrixConstantMem_15_io_data_4;
  wire       [254:0]  matrixConstantMem_16_io_data_0;
  wire       [254:0]  matrixConstantMem_16_io_data_1;
  wire       [254:0]  matrixConstantMem_16_io_data_2;
  wire       [254:0]  matrixConstantMem_16_io_data_3;
  wire       [254:0]  matrixConstantMem_16_io_data_4;
  wire       [254:0]  matrixConstantMem_16_io_data_5;
  wire       [254:0]  matrixConstantMem_16_io_data_6;
  wire       [254:0]  matrixConstantMem_16_io_data_7;
  wire       [254:0]  matrixConstantMem_16_io_data_8;
  wire       [254:0]  matrixConstantMem_17_io_data_0;
  wire       [254:0]  matrixConstantMem_17_io_data_1;
  wire       [254:0]  matrixConstantMem_17_io_data_2;
  wire       [254:0]  matrixConstantMem_17_io_data_3;
  wire       [254:0]  matrixConstantMem_17_io_data_4;
  wire       [254:0]  matrixConstantMem_17_io_data_5;
  wire       [254:0]  matrixConstantMem_17_io_data_6;
  wire       [254:0]  matrixConstantMem_17_io_data_7;
  wire       [254:0]  matrixConstantMem_17_io_data_8;
  wire       [254:0]  matrixConstantMem_17_io_data_9;
  wire       [254:0]  matrixConstantMem_17_io_data_10;
  wire       [254:0]  matrixConstantMem_17_io_data_11;
  wire       [254:0]  matrixConstantMem_18_io_data_0;
  wire       [254:0]  matrixConstantMem_18_io_data_1;
  wire       [254:0]  matrixConstantMem_18_io_data_2;
  wire       [254:0]  matrixConstantMem_19_io_data_0;
  wire       [254:0]  matrixConstantMem_19_io_data_1;
  wire       [254:0]  matrixConstantMem_19_io_data_2;
  wire       [254:0]  matrixConstantMem_19_io_data_3;
  wire       [254:0]  matrixConstantMem_19_io_data_4;
  wire       [254:0]  matrixConstantMem_20_io_data_0;
  wire       [254:0]  matrixConstantMem_20_io_data_1;
  wire       [254:0]  matrixConstantMem_20_io_data_2;
  wire       [254:0]  matrixConstantMem_20_io_data_3;
  wire       [254:0]  matrixConstantMem_20_io_data_4;
  wire       [254:0]  matrixConstantMem_20_io_data_5;
  wire       [254:0]  matrixConstantMem_20_io_data_6;
  wire       [254:0]  matrixConstantMem_20_io_data_7;
  wire       [254:0]  matrixConstantMem_20_io_data_8;
  wire       [254:0]  matrixConstantMem_21_io_data_0;
  wire       [254:0]  matrixConstantMem_21_io_data_1;
  wire       [254:0]  matrixConstantMem_21_io_data_2;
  wire       [254:0]  matrixConstantMem_21_io_data_3;
  wire       [254:0]  matrixConstantMem_21_io_data_4;
  wire       [254:0]  matrixConstantMem_21_io_data_5;
  wire       [254:0]  matrixConstantMem_21_io_data_6;
  wire       [254:0]  matrixConstantMem_21_io_data_7;
  wire       [254:0]  matrixConstantMem_21_io_data_8;
  wire       [254:0]  matrixConstantMem_21_io_data_9;
  wire       [254:0]  matrixConstantMem_21_io_data_10;
  wire       [254:0]  matrixConstantMem_21_io_data_11;
  wire       [254:0]  matrixConstantMem_22_io_data_0;
  wire       [254:0]  matrixConstantMem_22_io_data_1;
  wire       [254:0]  matrixConstantMem_22_io_data_2;
  wire       [254:0]  matrixConstantMem_22_io_data_3;
  wire       [254:0]  matrixConstantMem_22_io_data_4;
  wire       [254:0]  matrixConstantMem_23_io_data_0;
  wire       [254:0]  matrixConstantMem_23_io_data_1;
  wire       [254:0]  matrixConstantMem_23_io_data_2;
  wire       [254:0]  matrixConstantMem_23_io_data_3;
  wire       [254:0]  matrixConstantMem_23_io_data_4;
  wire       [254:0]  matrixConstantMem_23_io_data_5;
  wire       [254:0]  matrixConstantMem_23_io_data_6;
  wire       [254:0]  matrixConstantMem_23_io_data_7;
  wire       [254:0]  matrixConstantMem_23_io_data_8;
  wire       [254:0]  matrixConstantMem_24_io_data_0;
  wire       [254:0]  matrixConstantMem_24_io_data_1;
  wire       [254:0]  matrixConstantMem_24_io_data_2;
  wire       [254:0]  matrixConstantMem_24_io_data_3;
  wire       [254:0]  matrixConstantMem_24_io_data_4;
  wire       [254:0]  matrixConstantMem_24_io_data_5;
  wire       [254:0]  matrixConstantMem_24_io_data_6;
  wire       [254:0]  matrixConstantMem_24_io_data_7;
  wire       [254:0]  matrixConstantMem_24_io_data_8;
  wire       [254:0]  matrixConstantMem_25_io_data_0;
  wire       [254:0]  matrixConstantMem_25_io_data_1;
  wire       [254:0]  matrixConstantMem_25_io_data_2;
  wire       [254:0]  matrixConstantMem_25_io_data_3;
  wire       [254:0]  matrixConstantMem_25_io_data_4;
  wire       [254:0]  matrixConstantMem_25_io_data_5;
  wire       [254:0]  matrixConstantMem_25_io_data_6;
  wire       [254:0]  matrixConstantMem_25_io_data_7;
  wire       [254:0]  matrixConstantMem_25_io_data_8;
  wire       [254:0]  matrixConstantMem_25_io_data_9;
  wire       [254:0]  matrixConstantMem_25_io_data_10;
  wire       [254:0]  matrixConstantMem_25_io_data_11;
  wire       [254:0]  matrixConstantMem_26_io_data_0;
  wire       [254:0]  matrixConstantMem_26_io_data_1;
  wire       [254:0]  matrixConstantMem_26_io_data_2;
  wire       [254:0]  matrixConstantMem_26_io_data_3;
  wire       [254:0]  matrixConstantMem_26_io_data_4;
  wire       [254:0]  matrixConstantMem_26_io_data_5;
  wire       [254:0]  matrixConstantMem_26_io_data_6;
  wire       [254:0]  matrixConstantMem_26_io_data_7;
  wire       [254:0]  matrixConstantMem_26_io_data_8;
  wire       [254:0]  matrixConstantMem_27_io_data_0;
  wire       [254:0]  matrixConstantMem_27_io_data_1;
  wire       [254:0]  matrixConstantMem_27_io_data_2;
  wire       [254:0]  matrixConstantMem_27_io_data_3;
  wire       [254:0]  matrixConstantMem_27_io_data_4;
  wire       [254:0]  matrixConstantMem_27_io_data_5;
  wire       [254:0]  matrixConstantMem_27_io_data_6;
  wire       [254:0]  matrixConstantMem_27_io_data_7;
  wire       [254:0]  matrixConstantMem_27_io_data_8;
  wire       [254:0]  matrixConstantMem_27_io_data_9;
  wire       [254:0]  matrixConstantMem_27_io_data_10;
  wire       [254:0]  matrixConstantMem_27_io_data_11;
  wire       [764:0]  _zz_fullRound_mdsOutputs_0;
  wire       [1274:0] _zz_fullRound_mdsOutputs_1;
  wire       [2294:0] _zz_fullRound_mdsOutputs_2;
  wire       [3059:0] _zz_fullRound_mdsOutputs_3;
  wire       [254:0]  _zz_fullRound_mdsOutputs_3_1;
  wire       [254:0]  _zz_fullRound_mdsOutputs_3_2;
  reg        [3059:0] _zz_fullRound_mdsOutput_2;
  wire       [1:0]    _zz_fullRound_mdsOutput_3;
  wire       [764:0]  _zz_fullRound_preSparseOutputs_0;
  wire       [1274:0] _zz_fullRound_preSparseOutputs_1;
  wire       [2294:0] _zz_fullRound_preSparseOutputs_2;
  wire       [3059:0] _zz_fullRound_preSparseOutputs_3;
  wire       [254:0]  _zz_fullRound_preSparseOutputs_3_1;
  wire       [254:0]  _zz_fullRound_preSparseOutputs_3_2;
  reg        [3059:0] _zz_fullRound_preSparseOutput_2;
  wire       [1:0]    _zz_fullRound_preSparseOutput_3;
  wire       [254:0]  _zz_partialRound_sparseRowT12;
  wire       [254:0]  _zz_partialRound_sparseRowT12_1;
  wire       [254:0]  _zz_partialRound_sparseColT12;
  wire       [254:0]  _zz_partialRound_sparseColT12_1;
  wire       [1274:0] _zz_partialRound_sparseOutputs_0;
  wire       [2294:0] _zz_partialRound_sparseOutputs_1;
  reg        [3059:0] _zz_partialRound_output_2;
  wire       [1:0]    _zz_partialRound_output_3;
  reg        [3:0]    io_addr_stateSize_delay_1;
  reg        [3:0]    fullRound_sizeDelayed1;
  wire                fullRound_sizeSelect1_0;
  wire                fullRound_sizeSelect1_1;
  wire                fullRound_sizeSelect1_2;
  wire                fullRound_sizeSelect1_3;
  wire       [3059:0] fullRound_mdsOutputs_0;
  wire       [3059:0] fullRound_mdsOutputs_1;
  wire       [3059:0] fullRound_mdsOutputs_2;
  wire       [3059:0] fullRound_mdsOutputs_3;
  wire                _zz_fullRound_mdsOutput;
  wire                _zz_fullRound_mdsOutput_1;
  reg        [3059:0] fullRound_mdsOutput;
  reg        [3:0]    io_addr_stateSize_delay_1_1;
  reg        [3:0]    fullRound_sizeDelayed2;
  wire                fullRound_sizeSelect2_0;
  wire                fullRound_sizeSelect2_1;
  wire                fullRound_sizeSelect2_2;
  wire                fullRound_sizeSelect2_3;
  wire       [3059:0] fullRound_preSparseOutputs_0;
  wire       [3059:0] fullRound_preSparseOutputs_1;
  wire       [3059:0] fullRound_preSparseOutputs_2;
  wire       [3059:0] fullRound_preSparseOutputs_3;
  wire                _zz_fullRound_preSparseOutput;
  wire                _zz_fullRound_preSparseOutput_1;
  reg        [3059:0] fullRound_preSparseOutput;
  reg        [2:0]    io_addr_fullRound_delay_1;
  reg        [2:0]    io_addr_fullRound_delay_2;
  reg        [2:0]    fullRound_fullRoundDelayed;
  reg        [3059:0] fullRound_output;
  reg        [254:0]  partialRound_sparseMatT3_0;
  reg        [254:0]  partialRound_sparseMatT3_1;
  reg        [254:0]  partialRound_sparseMatT3_2;
  reg        [254:0]  partialRound_sparseMatT3_3;
  reg        [254:0]  partialRound_sparseMatT3_4;
  reg        [254:0]  partialRound_sparseMatT5_0;
  reg        [254:0]  partialRound_sparseMatT5_1;
  reg        [254:0]  partialRound_sparseMatT5_2;
  reg        [254:0]  partialRound_sparseMatT5_3;
  reg        [254:0]  partialRound_sparseMatT5_4;
  reg        [254:0]  partialRound_sparseMatT5_5;
  reg        [254:0]  partialRound_sparseMatT5_6;
  reg        [254:0]  partialRound_sparseMatT5_7;
  reg        [254:0]  partialRound_sparseMatT5_8;
  wire       [2294:0] partialRound_sparseRowT9;
  wire       [3059:0] partialRound_sparseRowT12;
  wire       [2294:0] partialRound_sparseColT9;
  wire       [3059:0] partialRound_sparseColT12;
  reg        [3:0]    io_addr_stateIndex_delay_1;
  reg        [3:0]    partialRound_indexDelayed1;
  reg        [3:0]    io_addr_stateIndex_delay_1_1;
  reg        [3:0]    partialRound_indexDelayed2;
  reg        [2294:0] partialRound_sparseMatT9;
  reg        [3059:0] partialRound_sparseMatT12;
  wire       [3059:0] partialRound_sparseOutputs_0;
  wire       [3059:0] partialRound_sparseOutputs_1;
  wire       [3059:0] partialRound_sparseOutputs_2;
  reg        [3:0]    io_addr_stateSize_delay_1_2;
  reg        [3:0]    io_addr_stateSize_delay_2;
  reg        [3:0]    partialRound_sizeDelayed;
  wire                partialRound_sizeSelect_0;
  wire                partialRound_sizeSelect_1;
  wire                partialRound_sizeSelect_2;
  wire                partialRound_sizeSelect_3;
  wire                _zz_partialRound_output;
  wire                _zz_partialRound_output_1;
  reg        [3059:0] partialRound_output;
  reg                 io_addr_isFull_delay_1;
  reg                 io_addr_isFull_delay_2;
  reg                 io_addr_isFull_delay_3;
  reg                 isFullDelayed;
  reg        [3059:0] _zz_io_data_0;

  assign _zz_fullRound_mdsOutputs_0 = {matrixConstantMem_14_io_data_2,{matrixConstantMem_14_io_data_1,matrixConstantMem_14_io_data_0}};
  assign _zz_fullRound_mdsOutputs_1 = {matrixConstantMem_15_io_data_4,{matrixConstantMem_15_io_data_3,{matrixConstantMem_15_io_data_2,{matrixConstantMem_15_io_data_1,matrixConstantMem_15_io_data_0}}}};
  assign _zz_fullRound_mdsOutputs_2 = {matrixConstantMem_16_io_data_8,{matrixConstantMem_16_io_data_7,{matrixConstantMem_16_io_data_6,{matrixConstantMem_16_io_data_5,{matrixConstantMem_16_io_data_4,{matrixConstantMem_16_io_data_3,{matrixConstantMem_16_io_data_2,{matrixConstantMem_16_io_data_1,matrixConstantMem_16_io_data_0}}}}}}}};
  assign _zz_fullRound_mdsOutputs_3 = {matrixConstantMem_17_io_data_11,{matrixConstantMem_17_io_data_10,{matrixConstantMem_17_io_data_9,{matrixConstantMem_17_io_data_8,{matrixConstantMem_17_io_data_7,{matrixConstantMem_17_io_data_6,{matrixConstantMem_17_io_data_5,{matrixConstantMem_17_io_data_4,{matrixConstantMem_17_io_data_3,{matrixConstantMem_17_io_data_2,{_zz_fullRound_mdsOutputs_3_1,_zz_fullRound_mdsOutputs_3_2}}}}}}}}}}};
  assign _zz_fullRound_preSparseOutputs_0 = {matrixConstantMem_18_io_data_2,{matrixConstantMem_18_io_data_1,matrixConstantMem_18_io_data_0}};
  assign _zz_fullRound_preSparseOutputs_1 = {matrixConstantMem_19_io_data_4,{matrixConstantMem_19_io_data_3,{matrixConstantMem_19_io_data_2,{matrixConstantMem_19_io_data_1,matrixConstantMem_19_io_data_0}}}};
  assign _zz_fullRound_preSparseOutputs_2 = {matrixConstantMem_20_io_data_8,{matrixConstantMem_20_io_data_7,{matrixConstantMem_20_io_data_6,{matrixConstantMem_20_io_data_5,{matrixConstantMem_20_io_data_4,{matrixConstantMem_20_io_data_3,{matrixConstantMem_20_io_data_2,{matrixConstantMem_20_io_data_1,matrixConstantMem_20_io_data_0}}}}}}}};
  assign _zz_fullRound_preSparseOutputs_3 = {matrixConstantMem_21_io_data_11,{matrixConstantMem_21_io_data_10,{matrixConstantMem_21_io_data_9,{matrixConstantMem_21_io_data_8,{matrixConstantMem_21_io_data_7,{matrixConstantMem_21_io_data_6,{matrixConstantMem_21_io_data_5,{matrixConstantMem_21_io_data_4,{matrixConstantMem_21_io_data_3,{matrixConstantMem_21_io_data_2,{_zz_fullRound_preSparseOutputs_3_1,_zz_fullRound_preSparseOutputs_3_2}}}}}}}}}}};
  assign _zz_partialRound_sparseOutputs_0 = {partialRound_sparseMatT3_4,{partialRound_sparseMatT3_3,{partialRound_sparseMatT3_2,{partialRound_sparseMatT3_1,partialRound_sparseMatT3_0}}}};
  assign _zz_partialRound_sparseOutputs_1 = {partialRound_sparseMatT5_8,{partialRound_sparseMatT5_7,{partialRound_sparseMatT5_6,{partialRound_sparseMatT5_5,{partialRound_sparseMatT5_4,{partialRound_sparseMatT5_3,{partialRound_sparseMatT5_2,{partialRound_sparseMatT5_1,partialRound_sparseMatT5_0}}}}}}}};
  assign _zz_fullRound_mdsOutput_3 = {_zz_fullRound_mdsOutput_1,_zz_fullRound_mdsOutput};
  assign _zz_fullRound_preSparseOutput_3 = {_zz_fullRound_preSparseOutput_1,_zz_fullRound_preSparseOutput};
  assign _zz_partialRound_output_3 = {_zz_partialRound_output_1,_zz_partialRound_output};
  assign _zz_fullRound_mdsOutputs_3_1 = matrixConstantMem_17_io_data_1;
  assign _zz_fullRound_mdsOutputs_3_2 = matrixConstantMem_17_io_data_0;
  assign _zz_fullRound_preSparseOutputs_3_1 = matrixConstantMem_21_io_data_1;
  assign _zz_fullRound_preSparseOutputs_3_2 = matrixConstantMem_21_io_data_0;
  assign _zz_partialRound_sparseRowT12 = matrixConstantMem_25_io_data_1;
  assign _zz_partialRound_sparseRowT12_1 = matrixConstantMem_25_io_data_0;
  assign _zz_partialRound_sparseColT12 = matrixConstantMem_27_io_data_1;
  assign _zz_partialRound_sparseColT12_1 = matrixConstantMem_27_io_data_0;
  MatrixConstantMem matrixConstantMem_14 (
    .io_data_0    (matrixConstantMem_14_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_14_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_14_io_data_2[254:0]  ), //o
    .io_addr      (matrixConstantMem_14_io_addr[1:0]      ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_1 matrixConstantMem_15 (
    .io_data_0    (matrixConstantMem_15_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_15_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_15_io_data_2[254:0]  ), //o
    .io_data_3    (matrixConstantMem_15_io_data_3[254:0]  ), //o
    .io_data_4    (matrixConstantMem_15_io_data_4[254:0]  ), //o
    .io_addr      (matrixConstantMem_15_io_addr[2:0]      ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_2 matrixConstantMem_16 (
    .io_data_0    (matrixConstantMem_16_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_16_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_16_io_data_2[254:0]  ), //o
    .io_data_3    (matrixConstantMem_16_io_data_3[254:0]  ), //o
    .io_data_4    (matrixConstantMem_16_io_data_4[254:0]  ), //o
    .io_data_5    (matrixConstantMem_16_io_data_5[254:0]  ), //o
    .io_data_6    (matrixConstantMem_16_io_data_6[254:0]  ), //o
    .io_data_7    (matrixConstantMem_16_io_data_7[254:0]  ), //o
    .io_data_8    (matrixConstantMem_16_io_data_8[254:0]  ), //o
    .io_addr      (io_addr_stateIndex[3:0]                ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_3 matrixConstantMem_17 (
    .io_data_0     (matrixConstantMem_17_io_data_0[254:0]   ), //o
    .io_data_1     (matrixConstantMem_17_io_data_1[254:0]   ), //o
    .io_data_2     (matrixConstantMem_17_io_data_2[254:0]   ), //o
    .io_data_3     (matrixConstantMem_17_io_data_3[254:0]   ), //o
    .io_data_4     (matrixConstantMem_17_io_data_4[254:0]   ), //o
    .io_data_5     (matrixConstantMem_17_io_data_5[254:0]   ), //o
    .io_data_6     (matrixConstantMem_17_io_data_6[254:0]   ), //o
    .io_data_7     (matrixConstantMem_17_io_data_7[254:0]   ), //o
    .io_data_8     (matrixConstantMem_17_io_data_8[254:0]   ), //o
    .io_data_9     (matrixConstantMem_17_io_data_9[254:0]   ), //o
    .io_data_10    (matrixConstantMem_17_io_data_10[254:0]  ), //o
    .io_data_11    (matrixConstantMem_17_io_data_11[254:0]  ), //o
    .io_addr       (io_addr_stateIndex[3:0]                 ), //i
    .clk           (clk                                     ), //i
    .resetn        (resetn                                  )  //i
  );
  MatrixConstantMem_4 matrixConstantMem_18 (
    .io_data_0    (matrixConstantMem_18_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_18_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_18_io_data_2[254:0]  ), //o
    .io_addr      (matrixConstantMem_18_io_addr[1:0]      ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_5 matrixConstantMem_19 (
    .io_data_0    (matrixConstantMem_19_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_19_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_19_io_data_2[254:0]  ), //o
    .io_data_3    (matrixConstantMem_19_io_data_3[254:0]  ), //o
    .io_data_4    (matrixConstantMem_19_io_data_4[254:0]  ), //o
    .io_addr      (matrixConstantMem_19_io_addr[2:0]      ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_6 matrixConstantMem_20 (
    .io_data_0    (matrixConstantMem_20_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_20_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_20_io_data_2[254:0]  ), //o
    .io_data_3    (matrixConstantMem_20_io_data_3[254:0]  ), //o
    .io_data_4    (matrixConstantMem_20_io_data_4[254:0]  ), //o
    .io_data_5    (matrixConstantMem_20_io_data_5[254:0]  ), //o
    .io_data_6    (matrixConstantMem_20_io_data_6[254:0]  ), //o
    .io_data_7    (matrixConstantMem_20_io_data_7[254:0]  ), //o
    .io_data_8    (matrixConstantMem_20_io_data_8[254:0]  ), //o
    .io_addr      (io_addr_stateIndex[3:0]                ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_7 matrixConstantMem_21 (
    .io_data_0     (matrixConstantMem_21_io_data_0[254:0]   ), //o
    .io_data_1     (matrixConstantMem_21_io_data_1[254:0]   ), //o
    .io_data_2     (matrixConstantMem_21_io_data_2[254:0]   ), //o
    .io_data_3     (matrixConstantMem_21_io_data_3[254:0]   ), //o
    .io_data_4     (matrixConstantMem_21_io_data_4[254:0]   ), //o
    .io_data_5     (matrixConstantMem_21_io_data_5[254:0]   ), //o
    .io_data_6     (matrixConstantMem_21_io_data_6[254:0]   ), //o
    .io_data_7     (matrixConstantMem_21_io_data_7[254:0]   ), //o
    .io_data_8     (matrixConstantMem_21_io_data_8[254:0]   ), //o
    .io_data_9     (matrixConstantMem_21_io_data_9[254:0]   ), //o
    .io_data_10    (matrixConstantMem_21_io_data_10[254:0]  ), //o
    .io_data_11    (matrixConstantMem_21_io_data_11[254:0]  ), //o
    .io_addr       (io_addr_stateIndex[3:0]                 ), //i
    .clk           (clk                                     ), //i
    .resetn        (resetn                                  )  //i
  );
  MatrixConstantMem_8 matrixConstantMem_22 (
    .io_data_0    (matrixConstantMem_22_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_22_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_22_io_data_2[254:0]  ), //o
    .io_data_3    (matrixConstantMem_22_io_data_3[254:0]  ), //o
    .io_data_4    (matrixConstantMem_22_io_data_4[254:0]  ), //o
    .io_addr      (io_addr_partialRound[5:0]              ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_9 matrixConstantMem_23 (
    .io_data_0    (matrixConstantMem_23_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_23_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_23_io_data_2[254:0]  ), //o
    .io_data_3    (matrixConstantMem_23_io_data_3[254:0]  ), //o
    .io_data_4    (matrixConstantMem_23_io_data_4[254:0]  ), //o
    .io_data_5    (matrixConstantMem_23_io_data_5[254:0]  ), //o
    .io_data_6    (matrixConstantMem_23_io_data_6[254:0]  ), //o
    .io_data_7    (matrixConstantMem_23_io_data_7[254:0]  ), //o
    .io_data_8    (matrixConstantMem_23_io_data_8[254:0]  ), //o
    .io_addr      (io_addr_partialRound[5:0]              ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_10 matrixConstantMem_24 (
    .io_data_0    (matrixConstantMem_24_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_24_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_24_io_data_2[254:0]  ), //o
    .io_data_3    (matrixConstantMem_24_io_data_3[254:0]  ), //o
    .io_data_4    (matrixConstantMem_24_io_data_4[254:0]  ), //o
    .io_data_5    (matrixConstantMem_24_io_data_5[254:0]  ), //o
    .io_data_6    (matrixConstantMem_24_io_data_6[254:0]  ), //o
    .io_data_7    (matrixConstantMem_24_io_data_7[254:0]  ), //o
    .io_data_8    (matrixConstantMem_24_io_data_8[254:0]  ), //o
    .io_addr      (io_addr_partialRound[5:0]              ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_11 matrixConstantMem_25 (
    .io_data_0     (matrixConstantMem_25_io_data_0[254:0]   ), //o
    .io_data_1     (matrixConstantMem_25_io_data_1[254:0]   ), //o
    .io_data_2     (matrixConstantMem_25_io_data_2[254:0]   ), //o
    .io_data_3     (matrixConstantMem_25_io_data_3[254:0]   ), //o
    .io_data_4     (matrixConstantMem_25_io_data_4[254:0]   ), //o
    .io_data_5     (matrixConstantMem_25_io_data_5[254:0]   ), //o
    .io_data_6     (matrixConstantMem_25_io_data_6[254:0]   ), //o
    .io_data_7     (matrixConstantMem_25_io_data_7[254:0]   ), //o
    .io_data_8     (matrixConstantMem_25_io_data_8[254:0]   ), //o
    .io_data_9     (matrixConstantMem_25_io_data_9[254:0]   ), //o
    .io_data_10    (matrixConstantMem_25_io_data_10[254:0]  ), //o
    .io_data_11    (matrixConstantMem_25_io_data_11[254:0]  ), //o
    .io_addr       (io_addr_partialRound[5:0]               ), //i
    .clk           (clk                                     ), //i
    .resetn        (resetn                                  )  //i
  );
  MatrixConstantMem_12 matrixConstantMem_26 (
    .io_data_0    (matrixConstantMem_26_io_data_0[254:0]  ), //o
    .io_data_1    (matrixConstantMem_26_io_data_1[254:0]  ), //o
    .io_data_2    (matrixConstantMem_26_io_data_2[254:0]  ), //o
    .io_data_3    (matrixConstantMem_26_io_data_3[254:0]  ), //o
    .io_data_4    (matrixConstantMem_26_io_data_4[254:0]  ), //o
    .io_data_5    (matrixConstantMem_26_io_data_5[254:0]  ), //o
    .io_data_6    (matrixConstantMem_26_io_data_6[254:0]  ), //o
    .io_data_7    (matrixConstantMem_26_io_data_7[254:0]  ), //o
    .io_data_8    (matrixConstantMem_26_io_data_8[254:0]  ), //o
    .io_addr      (io_addr_partialRound[5:0]              ), //i
    .clk          (clk                                    ), //i
    .resetn       (resetn                                 )  //i
  );
  MatrixConstantMem_13 matrixConstantMem_27 (
    .io_data_0     (matrixConstantMem_27_io_data_0[254:0]   ), //o
    .io_data_1     (matrixConstantMem_27_io_data_1[254:0]   ), //o
    .io_data_2     (matrixConstantMem_27_io_data_2[254:0]   ), //o
    .io_data_3     (matrixConstantMem_27_io_data_3[254:0]   ), //o
    .io_data_4     (matrixConstantMem_27_io_data_4[254:0]   ), //o
    .io_data_5     (matrixConstantMem_27_io_data_5[254:0]   ), //o
    .io_data_6     (matrixConstantMem_27_io_data_6[254:0]   ), //o
    .io_data_7     (matrixConstantMem_27_io_data_7[254:0]   ), //o
    .io_data_8     (matrixConstantMem_27_io_data_8[254:0]   ), //o
    .io_data_9     (matrixConstantMem_27_io_data_9[254:0]   ), //o
    .io_data_10    (matrixConstantMem_27_io_data_10[254:0]  ), //o
    .io_data_11    (matrixConstantMem_27_io_data_11[254:0]  ), //o
    .io_addr       (io_addr_partialRound[5:0]               ), //i
    .clk           (clk                                     ), //i
    .resetn        (resetn                                  )  //i
  );
  always @(*) begin
    case(_zz_fullRound_mdsOutput_3)
      2'b00 : _zz_fullRound_mdsOutput_2 = fullRound_mdsOutputs_0;
      2'b01 : _zz_fullRound_mdsOutput_2 = fullRound_mdsOutputs_1;
      2'b10 : _zz_fullRound_mdsOutput_2 = fullRound_mdsOutputs_2;
      default : _zz_fullRound_mdsOutput_2 = fullRound_mdsOutputs_3;
    endcase
  end

  always @(*) begin
    case(_zz_fullRound_preSparseOutput_3)
      2'b00 : _zz_fullRound_preSparseOutput_2 = fullRound_preSparseOutputs_0;
      2'b01 : _zz_fullRound_preSparseOutput_2 = fullRound_preSparseOutputs_1;
      2'b10 : _zz_fullRound_preSparseOutput_2 = fullRound_preSparseOutputs_2;
      default : _zz_fullRound_preSparseOutput_2 = fullRound_preSparseOutputs_3;
    endcase
  end

  always @(*) begin
    case(_zz_partialRound_output_3)
      2'b00 : _zz_partialRound_output_2 = partialRound_sparseOutputs_0;
      2'b01 : _zz_partialRound_output_2 = partialRound_sparseOutputs_1;
      2'b10 : _zz_partialRound_output_2 = partialRound_sparseOutputs_2;
      default : _zz_partialRound_output_2 = partialRound_sparseMatT12;
    endcase
  end

  assign fullRound_sizeSelect1_0 = (4'b0011 == fullRound_sizeDelayed1);
  assign fullRound_sizeSelect1_1 = (4'b0101 == fullRound_sizeDelayed1);
  assign fullRound_sizeSelect1_2 = (4'b1001 == fullRound_sizeDelayed1);
  assign fullRound_sizeSelect1_3 = (4'b1100 == fullRound_sizeDelayed1);
  assign matrixConstantMem_14_io_addr = io_addr_stateIndex[1:0];
  assign fullRound_mdsOutputs_0 = {2295'd0, _zz_fullRound_mdsOutputs_0};
  assign matrixConstantMem_15_io_addr = io_addr_stateIndex[2:0];
  assign fullRound_mdsOutputs_1 = {1785'd0, _zz_fullRound_mdsOutputs_1};
  assign fullRound_mdsOutputs_2 = {765'd0, _zz_fullRound_mdsOutputs_2};
  assign fullRound_mdsOutputs_3 = _zz_fullRound_mdsOutputs_3;
  assign _zz_fullRound_mdsOutput = (fullRound_sizeSelect1_1 || fullRound_sizeSelect1_3);
  assign _zz_fullRound_mdsOutput_1 = (fullRound_sizeSelect1_2 || fullRound_sizeSelect1_3);
  assign fullRound_sizeSelect2_0 = (4'b0011 == fullRound_sizeDelayed2);
  assign fullRound_sizeSelect2_1 = (4'b0101 == fullRound_sizeDelayed2);
  assign fullRound_sizeSelect2_2 = (4'b1001 == fullRound_sizeDelayed2);
  assign fullRound_sizeSelect2_3 = (4'b1100 == fullRound_sizeDelayed2);
  assign matrixConstantMem_18_io_addr = io_addr_stateIndex[1:0];
  assign fullRound_preSparseOutputs_0 = {2295'd0, _zz_fullRound_preSparseOutputs_0};
  assign matrixConstantMem_19_io_addr = io_addr_stateIndex[2:0];
  assign fullRound_preSparseOutputs_1 = {1785'd0, _zz_fullRound_preSparseOutputs_1};
  assign fullRound_preSparseOutputs_2 = {765'd0, _zz_fullRound_preSparseOutputs_2};
  assign fullRound_preSparseOutputs_3 = _zz_fullRound_preSparseOutputs_3;
  assign _zz_fullRound_preSparseOutput = (fullRound_sizeSelect2_1 || fullRound_sizeSelect2_3);
  assign _zz_fullRound_preSparseOutput_1 = (fullRound_sizeSelect2_2 || fullRound_sizeSelect2_3);
  assign partialRound_sparseRowT9 = {matrixConstantMem_24_io_data_8,{matrixConstantMem_24_io_data_7,{matrixConstantMem_24_io_data_6,{matrixConstantMem_24_io_data_5,{matrixConstantMem_24_io_data_4,{matrixConstantMem_24_io_data_3,{matrixConstantMem_24_io_data_2,{matrixConstantMem_24_io_data_1,matrixConstantMem_24_io_data_0}}}}}}}};
  assign partialRound_sparseRowT12 = {matrixConstantMem_25_io_data_11,{matrixConstantMem_25_io_data_10,{matrixConstantMem_25_io_data_9,{matrixConstantMem_25_io_data_8,{matrixConstantMem_25_io_data_7,{matrixConstantMem_25_io_data_6,{matrixConstantMem_25_io_data_5,{matrixConstantMem_25_io_data_4,{matrixConstantMem_25_io_data_3,{matrixConstantMem_25_io_data_2,{_zz_partialRound_sparseRowT12,_zz_partialRound_sparseRowT12_1}}}}}}}}}}};
  assign partialRound_sparseColT9 = {matrixConstantMem_26_io_data_8,{matrixConstantMem_26_io_data_7,{matrixConstantMem_26_io_data_6,{matrixConstantMem_26_io_data_5,{matrixConstantMem_26_io_data_4,{matrixConstantMem_26_io_data_3,{matrixConstantMem_26_io_data_2,{matrixConstantMem_26_io_data_1,matrixConstantMem_26_io_data_0}}}}}}}};
  assign partialRound_sparseColT12 = {matrixConstantMem_27_io_data_11,{matrixConstantMem_27_io_data_10,{matrixConstantMem_27_io_data_9,{matrixConstantMem_27_io_data_8,{matrixConstantMem_27_io_data_7,{matrixConstantMem_27_io_data_6,{matrixConstantMem_27_io_data_5,{matrixConstantMem_27_io_data_4,{matrixConstantMem_27_io_data_3,{matrixConstantMem_27_io_data_2,{_zz_partialRound_sparseColT12,_zz_partialRound_sparseColT12_1}}}}}}}}}}};
  assign partialRound_sparseOutputs_0 = {1785'd0, _zz_partialRound_sparseOutputs_0};
  assign partialRound_sparseOutputs_1 = {765'd0, _zz_partialRound_sparseOutputs_1};
  assign partialRound_sparseOutputs_2 = {765'd0, partialRound_sparseMatT9};
  assign partialRound_sizeSelect_0 = (4'b0011 == partialRound_sizeDelayed);
  assign partialRound_sizeSelect_1 = (4'b0101 == partialRound_sizeDelayed);
  assign partialRound_sizeSelect_2 = (4'b1001 == partialRound_sizeDelayed);
  assign partialRound_sizeSelect_3 = (4'b1100 == partialRound_sizeDelayed);
  assign _zz_partialRound_output = (partialRound_sizeSelect_1 || partialRound_sizeSelect_3);
  assign _zz_partialRound_output_1 = (partialRound_sizeSelect_2 || partialRound_sizeSelect_3);
  assign io_data_0 = _zz_io_data_0[254 : 0];
  assign io_data_1 = _zz_io_data_0[509 : 255];
  assign io_data_2 = _zz_io_data_0[764 : 510];
  assign io_data_3 = _zz_io_data_0[1019 : 765];
  assign io_data_4 = _zz_io_data_0[1274 : 1020];
  assign io_data_5 = _zz_io_data_0[1529 : 1275];
  assign io_data_6 = _zz_io_data_0[1784 : 1530];
  assign io_data_7 = _zz_io_data_0[2039 : 1785];
  assign io_data_8 = _zz_io_data_0[2294 : 2040];
  assign io_data_9 = _zz_io_data_0[2549 : 2295];
  assign io_data_10 = _zz_io_data_0[2804 : 2550];
  assign io_data_11 = _zz_io_data_0[3059 : 2805];
  always @(posedge clk) begin
    io_addr_stateSize_delay_1 <= io_addr_stateSize;
    fullRound_sizeDelayed1 <= io_addr_stateSize_delay_1;
    fullRound_mdsOutput <= _zz_fullRound_mdsOutput_2;
    io_addr_stateSize_delay_1_1 <= io_addr_stateSize;
    fullRound_sizeDelayed2 <= io_addr_stateSize_delay_1_1;
    fullRound_preSparseOutput <= _zz_fullRound_preSparseOutput_2;
    io_addr_fullRound_delay_1 <= io_addr_fullRound;
    io_addr_fullRound_delay_2 <= io_addr_fullRound_delay_1;
    fullRound_fullRoundDelayed <= io_addr_fullRound_delay_2;
    fullRound_output <= ((fullRound_fullRoundDelayed == 3'b011) ? fullRound_preSparseOutput : fullRound_mdsOutput);
    partialRound_sparseMatT3_0 <= matrixConstantMem_22_io_data_0;
    partialRound_sparseMatT3_1 <= matrixConstantMem_22_io_data_1;
    partialRound_sparseMatT3_2 <= matrixConstantMem_22_io_data_2;
    partialRound_sparseMatT3_3 <= matrixConstantMem_22_io_data_3;
    partialRound_sparseMatT3_4 <= matrixConstantMem_22_io_data_4;
    partialRound_sparseMatT5_0 <= matrixConstantMem_23_io_data_0;
    partialRound_sparseMatT5_1 <= matrixConstantMem_23_io_data_1;
    partialRound_sparseMatT5_2 <= matrixConstantMem_23_io_data_2;
    partialRound_sparseMatT5_3 <= matrixConstantMem_23_io_data_3;
    partialRound_sparseMatT5_4 <= matrixConstantMem_23_io_data_4;
    partialRound_sparseMatT5_5 <= matrixConstantMem_23_io_data_5;
    partialRound_sparseMatT5_6 <= matrixConstantMem_23_io_data_6;
    partialRound_sparseMatT5_7 <= matrixConstantMem_23_io_data_7;
    partialRound_sparseMatT5_8 <= matrixConstantMem_23_io_data_8;
    io_addr_stateIndex_delay_1 <= io_addr_stateIndex;
    partialRound_indexDelayed1 <= io_addr_stateIndex_delay_1;
    io_addr_stateIndex_delay_1_1 <= io_addr_stateIndex;
    partialRound_indexDelayed2 <= io_addr_stateIndex_delay_1_1;
    partialRound_sparseMatT9 <= ((partialRound_indexDelayed1 == 4'b0000) ? partialRound_sparseRowT9 : partialRound_sparseColT9);
    partialRound_sparseMatT12 <= ((partialRound_indexDelayed2 == 4'b0000) ? partialRound_sparseRowT12 : partialRound_sparseColT12);
    io_addr_stateSize_delay_1_2 <= io_addr_stateSize;
    io_addr_stateSize_delay_2 <= io_addr_stateSize_delay_1_2;
    partialRound_sizeDelayed <= io_addr_stateSize_delay_2;
    partialRound_output <= _zz_partialRound_output_2;
    io_addr_isFull_delay_1 <= io_addr_isFull;
    io_addr_isFull_delay_2 <= io_addr_isFull_delay_1;
    io_addr_isFull_delay_3 <= io_addr_isFull_delay_2;
    isFullDelayed <= io_addr_isFull_delay_3;
    _zz_io_data_0 <= (isFullDelayed ? fullRound_output : partialRound_output);
  end


endmodule

//AdderIPFlow replaced by AdderIPFlow

module AdderIPFlow (
  input               io_input_valid,
  input      [254:0]  io_input_payload_op1,
  input      [254:0]  io_input_payload_op2,
  output              io_output_valid,
  output     [255:0]  io_output_payload_res,
  input               clk,
  input               resetn
);

  wire       [255:0]  simAdderIP_48_io_outputS;
  reg                 io_input_valid_delay_1;
  reg                 io_input_valid_delay_2;
  reg                 io_input_valid_delay_3;
  reg                 io_input_valid_delay_4;
  reg                 io_input_valid_delay_5;
  reg                 io_input_valid_delay_6;
  reg                 io_input_valid_delay_7;
  reg                 io_input_valid_delay_8;
  reg                 io_input_valid_delay_9;
  reg                 io_input_valid_delay_10;
  reg                 io_input_valid_delay_11;
  reg                 io_input_valid_delay_12;
  reg                 io_input_valid_delay_13;
  reg                 io_input_valid_delay_14;
  reg                 io_input_valid_delay_15;
  reg                 validDelayed;

  SimAdderIP_22 simAdderIP_48 (
    .io_inputA     (io_input_payload_op1[254:0]      ), //i
    .io_inputB     (io_input_payload_op2[254:0]      ), //i
    .io_outputS    (simAdderIP_48_io_outputS[255:0]  ), //o
    .clk           (clk                              ), //i
    .resetn        (resetn                           )  //i
  );
  assign io_output_valid = validDelayed;
  assign io_output_payload_res = simAdderIP_48_io_outputS;
  always @(posedge clk) begin
    if(!resetn) begin
      io_input_valid_delay_1 <= 1'b0;
      io_input_valid_delay_2 <= 1'b0;
      io_input_valid_delay_3 <= 1'b0;
      io_input_valid_delay_4 <= 1'b0;
      io_input_valid_delay_5 <= 1'b0;
      io_input_valid_delay_6 <= 1'b0;
      io_input_valid_delay_7 <= 1'b0;
      io_input_valid_delay_8 <= 1'b0;
      io_input_valid_delay_9 <= 1'b0;
      io_input_valid_delay_10 <= 1'b0;
      io_input_valid_delay_11 <= 1'b0;
      io_input_valid_delay_12 <= 1'b0;
      io_input_valid_delay_13 <= 1'b0;
      io_input_valid_delay_14 <= 1'b0;
      io_input_valid_delay_15 <= 1'b0;
      validDelayed <= 1'b0;
    end else begin
      io_input_valid_delay_1 <= io_input_valid;
      io_input_valid_delay_2 <= io_input_valid_delay_1;
      io_input_valid_delay_3 <= io_input_valid_delay_2;
      io_input_valid_delay_4 <= io_input_valid_delay_3;
      io_input_valid_delay_5 <= io_input_valid_delay_4;
      io_input_valid_delay_6 <= io_input_valid_delay_5;
      io_input_valid_delay_7 <= io_input_valid_delay_6;
      io_input_valid_delay_8 <= io_input_valid_delay_7;
      io_input_valid_delay_9 <= io_input_valid_delay_8;
      io_input_valid_delay_10 <= io_input_valid_delay_9;
      io_input_valid_delay_11 <= io_input_valid_delay_10;
      io_input_valid_delay_12 <= io_input_valid_delay_11;
      io_input_valid_delay_13 <= io_input_valid_delay_12;
      io_input_valid_delay_14 <= io_input_valid_delay_13;
      io_input_valid_delay_15 <= io_input_valid_delay_14;
      validDelayed <= io_input_valid_delay_15;
    end
  end


endmodule

module PartialRoundConstantMem (
  input      [3:0]    io_stateSize,
  input      [5:0]    io_partialRound,
  output     [254:0]  io_constant
);

  wire       [254:0]  _zz_constantsMem_0_port0;
  wire       [254:0]  _zz_constantsMem_1_port0;
  wire       [254:0]  _zz_constantsMem_2_port0;
  wire       [254:0]  _zz_constantsMem_3_port0;
  reg        [254:0]  _zz_io_constant_2;
  wire       [1:0]    _zz_io_constant_3;
  wire       [251:0]  initialContent_0_0;
  wire       [254:0]  initialContent_0_1;
  wire       [246:0]  initialContent_0_2;
  wire       [254:0]  initialContent_0_3;
  wire       [253:0]  initialContent_0_4;
  wire       [254:0]  initialContent_0_5;
  wire       [250:0]  initialContent_0_6;
  wire       [253:0]  initialContent_0_7;
  wire       [254:0]  initialContent_0_8;
  wire       [253:0]  initialContent_0_9;
  wire       [252:0]  initialContent_0_10;
  wire       [253:0]  initialContent_0_11;
  wire       [252:0]  initialContent_0_12;
  wire       [254:0]  initialContent_0_13;
  wire       [249:0]  initialContent_0_14;
  wire       [251:0]  initialContent_0_15;
  wire       [254:0]  initialContent_0_16;
  wire       [251:0]  initialContent_0_17;
  wire       [254:0]  initialContent_0_18;
  wire       [254:0]  initialContent_0_19;
  wire       [252:0]  initialContent_0_20;
  wire       [252:0]  initialContent_0_21;
  wire       [252:0]  initialContent_0_22;
  wire       [252:0]  initialContent_0_23;
  wire       [253:0]  initialContent_0_24;
  wire       [253:0]  initialContent_0_25;
  wire       [253:0]  initialContent_0_26;
  wire       [254:0]  initialContent_0_27;
  wire       [251:0]  initialContent_0_28;
  wire       [254:0]  initialContent_0_29;
  wire       [254:0]  initialContent_0_30;
  wire       [254:0]  initialContent_0_31;
  wire       [254:0]  initialContent_0_32;
  wire       [253:0]  initialContent_0_33;
  wire       [254:0]  initialContent_0_34;
  wire       [254:0]  initialContent_0_35;
  wire       [251:0]  initialContent_0_36;
  wire       [254:0]  initialContent_0_37;
  wire       [253:0]  initialContent_0_38;
  wire       [253:0]  initialContent_0_39;
  wire       [251:0]  initialContent_0_40;
  wire       [252:0]  initialContent_0_41;
  wire       [254:0]  initialContent_0_42;
  wire       [253:0]  initialContent_0_43;
  wire       [254:0]  initialContent_0_44;
  wire       [254:0]  initialContent_0_45;
  wire       [254:0]  initialContent_0_46;
  wire       [253:0]  initialContent_0_47;
  wire       [254:0]  initialContent_0_48;
  wire       [254:0]  initialContent_0_49;
  wire       [253:0]  initialContent_0_50;
  wire       [253:0]  initialContent_0_51;
  wire       [254:0]  initialContent_0_52;
  wire       [254:0]  initialContent_0_53;
  wire       [253:0]  initialContent_0_54;
  wire       [254:0]  initialContent_1_0;
  wire       [254:0]  initialContent_1_1;
  wire       [253:0]  initialContent_1_2;
  wire       [251:0]  initialContent_1_3;
  wire       [254:0]  initialContent_1_4;
  wire       [254:0]  initialContent_1_5;
  wire       [252:0]  initialContent_1_6;
  wire       [253:0]  initialContent_1_7;
  wire       [252:0]  initialContent_1_8;
  wire       [250:0]  initialContent_1_9;
  wire       [254:0]  initialContent_1_10;
  wire       [254:0]  initialContent_1_11;
  wire       [253:0]  initialContent_1_12;
  wire       [254:0]  initialContent_1_13;
  wire       [254:0]  initialContent_1_14;
  wire       [251:0]  initialContent_1_15;
  wire       [253:0]  initialContent_1_16;
  wire       [253:0]  initialContent_1_17;
  wire       [254:0]  initialContent_1_18;
  wire       [252:0]  initialContent_1_19;
  wire       [254:0]  initialContent_1_20;
  wire       [250:0]  initialContent_1_21;
  wire       [251:0]  initialContent_1_22;
  wire       [254:0]  initialContent_1_23;
  wire       [252:0]  initialContent_1_24;
  wire       [254:0]  initialContent_1_25;
  wire       [252:0]  initialContent_1_26;
  wire       [250:0]  initialContent_1_27;
  wire       [254:0]  initialContent_1_28;
  wire       [254:0]  initialContent_1_29;
  wire       [254:0]  initialContent_1_30;
  wire       [252:0]  initialContent_1_31;
  wire       [253:0]  initialContent_1_32;
  wire       [253:0]  initialContent_1_33;
  wire       [254:0]  initialContent_1_34;
  wire       [254:0]  initialContent_1_35;
  wire       [250:0]  initialContent_1_36;
  wire       [254:0]  initialContent_1_37;
  wire       [251:0]  initialContent_1_38;
  wire       [253:0]  initialContent_1_39;
  wire       [253:0]  initialContent_1_40;
  wire       [254:0]  initialContent_1_41;
  wire       [253:0]  initialContent_1_42;
  wire       [253:0]  initialContent_1_43;
  wire       [254:0]  initialContent_1_44;
  wire       [253:0]  initialContent_1_45;
  wire       [253:0]  initialContent_1_46;
  wire       [254:0]  initialContent_1_47;
  wire       [252:0]  initialContent_1_48;
  wire       [251:0]  initialContent_1_49;
  wire       [254:0]  initialContent_1_50;
  wire       [252:0]  initialContent_1_51;
  wire       [254:0]  initialContent_1_52;
  wire       [254:0]  initialContent_1_53;
  wire       [247:0]  initialContent_1_54;
  wire       [254:0]  initialContent_1_55;
  wire       [254:0]  initialContent_2_0;
  wire       [254:0]  initialContent_2_1;
  wire       [254:0]  initialContent_2_2;
  wire       [254:0]  initialContent_2_3;
  wire       [253:0]  initialContent_2_4;
  wire       [254:0]  initialContent_2_5;
  wire       [251:0]  initialContent_2_6;
  wire       [254:0]  initialContent_2_7;
  wire       [254:0]  initialContent_2_8;
  wire       [249:0]  initialContent_2_9;
  wire       [252:0]  initialContent_2_10;
  wire       [254:0]  initialContent_2_11;
  wire       [254:0]  initialContent_2_12;
  wire       [251:0]  initialContent_2_13;
  wire       [252:0]  initialContent_2_14;
  wire       [253:0]  initialContent_2_15;
  wire       [253:0]  initialContent_2_16;
  wire       [254:0]  initialContent_2_17;
  wire       [254:0]  initialContent_2_18;
  wire       [253:0]  initialContent_2_19;
  wire       [254:0]  initialContent_2_20;
  wire       [251:0]  initialContent_2_21;
  wire       [251:0]  initialContent_2_22;
  wire       [252:0]  initialContent_2_23;
  wire       [254:0]  initialContent_2_24;
  wire       [254:0]  initialContent_2_25;
  wire       [254:0]  initialContent_2_26;
  wire       [254:0]  initialContent_2_27;
  wire       [254:0]  initialContent_2_28;
  wire       [253:0]  initialContent_2_29;
  wire       [254:0]  initialContent_2_30;
  wire       [253:0]  initialContent_2_31;
  wire       [251:0]  initialContent_2_32;
  wire       [254:0]  initialContent_2_33;
  wire       [250:0]  initialContent_2_34;
  wire       [253:0]  initialContent_2_35;
  wire       [254:0]  initialContent_2_36;
  wire       [253:0]  initialContent_2_37;
  wire       [253:0]  initialContent_2_38;
  wire       [254:0]  initialContent_2_39;
  wire       [252:0]  initialContent_2_40;
  wire       [252:0]  initialContent_2_41;
  wire       [253:0]  initialContent_2_42;
  wire       [254:0]  initialContent_2_43;
  wire       [254:0]  initialContent_2_44;
  wire       [254:0]  initialContent_2_45;
  wire       [251:0]  initialContent_2_46;
  wire       [254:0]  initialContent_2_47;
  wire       [253:0]  initialContent_2_48;
  wire       [254:0]  initialContent_2_49;
  wire       [253:0]  initialContent_2_50;
  wire       [251:0]  initialContent_2_51;
  wire       [253:0]  initialContent_2_52;
  wire       [254:0]  initialContent_2_53;
  wire       [254:0]  initialContent_2_54;
  wire       [253:0]  initialContent_2_55;
  wire       [254:0]  initialContent_2_56;
  wire       [254:0]  initialContent_3_0;
  wire       [253:0]  initialContent_3_1;
  wire       [253:0]  initialContent_3_2;
  wire       [253:0]  initialContent_3_3;
  wire       [253:0]  initialContent_3_4;
  wire       [252:0]  initialContent_3_5;
  wire       [254:0]  initialContent_3_6;
  wire       [254:0]  initialContent_3_7;
  wire       [254:0]  initialContent_3_8;
  wire       [254:0]  initialContent_3_9;
  wire       [254:0]  initialContent_3_10;
  wire       [249:0]  initialContent_3_11;
  wire       [252:0]  initialContent_3_12;
  wire       [254:0]  initialContent_3_13;
  wire       [251:0]  initialContent_3_14;
  wire       [248:0]  initialContent_3_15;
  wire       [254:0]  initialContent_3_16;
  wire       [253:0]  initialContent_3_17;
  wire       [253:0]  initialContent_3_18;
  wire       [252:0]  initialContent_3_19;
  wire       [251:0]  initialContent_3_20;
  wire       [254:0]  initialContent_3_21;
  wire       [254:0]  initialContent_3_22;
  wire       [254:0]  initialContent_3_23;
  wire       [253:0]  initialContent_3_24;
  wire       [254:0]  initialContent_3_25;
  wire       [254:0]  initialContent_3_26;
  wire       [254:0]  initialContent_3_27;
  wire       [253:0]  initialContent_3_28;
  wire       [254:0]  initialContent_3_29;
  wire       [253:0]  initialContent_3_30;
  wire       [254:0]  initialContent_3_31;
  wire       [253:0]  initialContent_3_32;
  wire       [253:0]  initialContent_3_33;
  wire       [254:0]  initialContent_3_34;
  wire       [253:0]  initialContent_3_35;
  wire       [252:0]  initialContent_3_36;
  wire       [254:0]  initialContent_3_37;
  wire       [254:0]  initialContent_3_38;
  wire       [254:0]  initialContent_3_39;
  wire       [254:0]  initialContent_3_40;
  wire       [253:0]  initialContent_3_41;
  wire       [254:0]  initialContent_3_42;
  wire       [252:0]  initialContent_3_43;
  wire       [254:0]  initialContent_3_44;
  wire       [252:0]  initialContent_3_45;
  wire       [253:0]  initialContent_3_46;
  wire       [249:0]  initialContent_3_47;
  wire       [254:0]  initialContent_3_48;
  wire       [253:0]  initialContent_3_49;
  wire       [253:0]  initialContent_3_50;
  wire       [254:0]  initialContent_3_51;
  wire       [249:0]  initialContent_3_52;
  wire       [253:0]  initialContent_3_53;
  wire       [254:0]  initialContent_3_54;
  wire       [252:0]  initialContent_3_55;
  wire       [251:0]  initialContent_3_56;
  wire       [5:0]    _zz_memOutputs_0;
  wire       [254:0]  memOutputs_0;
  wire       [5:0]    _zz_memOutputs_1;
  wire       [254:0]  memOutputs_1;
  wire       [5:0]    _zz_memOutputs_2;
  wire       [254:0]  memOutputs_2;
  wire       [5:0]    _zz_memOutputs_3;
  wire       [254:0]  memOutputs_3;
  wire                select_0;
  wire                select_1;
  wire                select_2;
  wire                select_3;
  wire                _zz_io_constant;
  wire                _zz_io_constant_1;
  (* ram_style = "distributed" *) reg [254:0] constantsMem_0 [0:54];
  (* ram_style = "distributed" *) reg [254:0] constantsMem_1 [0:55];
  (* ram_style = "distributed" *) reg [254:0] constantsMem_2 [0:56];
  (* ram_style = "distributed" *) reg [254:0] constantsMem_3 [0:56];

  assign _zz_io_constant_3 = {_zz_io_constant_1,_zz_io_constant};
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_partialRoundConstantMem_1_constantsMem_0.bin",constantsMem_0);
  end
  assign _zz_constantsMem_0_port0 = constantsMem_0[_zz_memOutputs_0];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_partialRoundConstantMem_1_constantsMem_1.bin",constantsMem_1);
  end
  assign _zz_constantsMem_1_port0 = constantsMem_1[_zz_memOutputs_1];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_partialRoundConstantMem_1_constantsMem_2.bin",constantsMem_2);
  end
  assign _zz_constantsMem_2_port0 = constantsMem_2[_zz_memOutputs_2];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_partialRoundConstantMem_1_constantsMem_3.bin",constantsMem_3);
  end
  assign _zz_constantsMem_3_port0 = constantsMem_3[_zz_memOutputs_3];
  always @(*) begin
    case(_zz_io_constant_3)
      2'b00 : _zz_io_constant_2 = memOutputs_0;
      2'b01 : _zz_io_constant_2 = memOutputs_1;
      2'b10 : _zz_io_constant_2 = memOutputs_2;
      default : _zz_io_constant_2 = memOutputs_3;
    endcase
  end

  assign initialContent_0_0 = 252'h955a904fbfcb90fbc5defc5c7e2c54155cd6d72beae79db3270aeb7b2d94f2c;
  assign initialContent_0_1 = 255'h48f5beee5b2bdab502cc5b8c2ed81366933e432e83f45112b3c600d678069561;
  assign initialContent_0_2 = 247'h5e4d218e2cbf432276a71b1172e3e870bc72581a32e4cb320fbab29868befe;
  assign initialContent_0_3 = 255'h40786413d77419f01c1f4b55932d717d6dd60a3567f47a00f192f40a6de7145b;
  assign initialContent_0_4 = 254'h21053c08db804c9ed0850bbd5200bc4cb4e51b9ccf99a93b97568646c2f5a9f2;
  assign initialContent_0_5 = 255'h696dcdc86c83f99b7ab110a0363b3e3be6ba21155fba71a5e33c6a07000694da;
  assign initialContent_0_6 = 251'h79e5780173271b97ad33f244e58cf742033f30121bb07a768eb1660c943a8cb;
  assign initialContent_0_7 = 254'h2ae60b92394ee0af5bcf1b75334c09b42b141c597f98f6ccee459235b5e7089d;
  assign initialContent_0_8 = 255'h6ca1fe4acfb19a5bc717c9dba926361ae42dc45ce97502696bd4c7dc43dd73e2;
  assign initialContent_0_9 = 254'h3213b3fa85b5ecda7f7a545e795072a3ccb959e291cedf0a44b4c0f3c3b3e539;
  assign initialContent_0_10 = 253'h1ae21be5ce235400a519d058a42cba01dbcfa358bd9f184609798ec6a14d217a;
  assign initialContent_0_11 = 254'h2e0d7726f80fb61131c55f1c9716450bc693731219d48bfc23c750fa2d8d28a1;
  assign initialContent_0_12 = 253'h181b74f358c9e32cfd1f921edd308e6a7fdb7c134231a08a820560707ea741ad;
  assign initialContent_0_13 = 255'h60719327c018006c11add949b16ac05bdda8bbd024ca707d8f3dbd3561c84ee9;
  assign initialContent_0_14 = 250'h2a278c8df95f69d8a3e968c60b5272cc0618b2b67efc17f938c3b7c49c9d2a8;
  assign initialContent_0_15 = 252'hb4820817e915168634f8adaf951f93cfd2d51996c9090050c3e1c16537432e2;
  assign initialContent_0_16 = 255'h463dfbe202dd6fe926bd3e67dc0e0819ce260112368084f23447e04fb812d49a;
  assign initialContent_0_17 = 252'h8e354ca57e78ee68ab9521c305d8a0c34ccdbded694b9e1f87ee0d9e01aca4e;
  assign initialContent_0_18 = 255'h5f0fe54b3ba4666e107322d50c08af509f062c46cf86264edb4ba5221412ae94;
  assign initialContent_0_19 = 255'h6414ea3cce47f294c4ef7587a070b7fd577faf359c64f44190e5c7c5d11c0582;
  assign initialContent_0_20 = 253'h17f8d17b6f8a1a89bd02f67dc8be4f78356d12a3769c6d277127a0c3bb978d48;
  assign initialContent_0_21 = 253'h1b64219f9c0bbcda51ca7f66c7ce4359dc57157a2831146ca3ca2266320004b6;
  assign initialContent_0_22 = 253'h10c0b3db7560da95d001063291d42a2715ea388788faf42d2832105acaaf128c;
  assign initialContent_0_23 = 253'h197aaac31652ed74fb001ff6203bb5eae7ca7c5069b7fb11514dd01cda3bcfba;
  assign initialContent_0_24 = 254'h38db32f5eea5fa8059d6e14534b4a7d7c06a3c6b4b93b7ba0519c9abb7a6fa36;
  assign initialContent_0_25 = 254'h34486da53591db38d19727c8ed2d7d4ea3077f27b533b7e629f26572656a8b08;
  assign initialContent_0_26 = 254'h24a138017e08c10f603a428b172054211ea417fea26618521c0aa85514af00e3;
  assign initialContent_0_27 = 255'h4d307087ecc872c0d08c5e961a8fa958cb35bb1067242fb2a91687266d874347;
  assign initialContent_0_28 = 252'hdcf58841afa7f5546ba57793eb05ac1e6b6de63628554a45f1bb36c5e2a1827;
  assign initialContent_0_29 = 255'h55fa9a0dba68e0a58207cddb42ff6a5d85a05677fe2b8bc2a12f1024bf6c96e5;
  assign initialContent_0_30 = 255'h7326ff2dcf3c878ecfd6d20491fa3d963cfe5e7bcd013806ec6556cef7c925e1;
  assign initialContent_0_31 = 255'h5e60fe3c2bea6ca8efadc4b05e47876297e63a714f2e13f62937f7282c3a87dd;
  assign initialContent_0_32 = 255'h5c5f684f78c673743fcdfbef6a307d255de584513584aa761430fdc74d7b0ea3;
  assign initialContent_0_33 = 254'h21639f6b8a8979ed5f546bb8cd0f7b9bbaf33d3e65fd6a3518ddae6fb61d4dd5;
  assign initialContent_0_34 = 255'h681903730747e00f2cc1958eddb0ebb0bd9a38a8468890a40e91f250640324b4;
  assign initialContent_0_35 = 255'h4fd7686552c2706f5b6007b1155fc62ae6c0664cc9630d2c81e3c47f0fdb7918;
  assign initialContent_0_36 = 252'hc36c60cf0bb29cd26509015a7e00681e698b79349aba3ff5e49924ff37d1138;
  assign initialContent_0_37 = 255'h487a6367936f46b7a017c850f166c30b6841bd1e96446da4d6dda0af276a82ad;
  assign initialContent_0_38 = 254'h36fb0be312dd473fc81b749586ecc089a940ce532efb5c1f92ed3f92ffdfee95;
  assign initialContent_0_39 = 254'h37963b1d7716c1fdde3829102d8f7a93ea75b4747573c9cee5a8514792db59ef;
  assign initialContent_0_40 = 252'h82045aa3c764242d6201cd77ddb4c9c03a217bba94eaa40a051faf3ebfe3cca;
  assign initialContent_0_41 = 253'h118af6e575fa8a991e7cbbd42ce8d65132d0d4ec3ee48d7ec6e45434ce32ee3f;
  assign initialContent_0_42 = 255'h5d08bf87451c7afff5ea4367a7fef5fc820d9f82c14c1f7045e734f865d9619e;
  assign initialContent_0_43 = 254'h214218ce6c8049edea3ee22f6aaf01892cb586efdd0591f73c3f44281fe9bf6b;
  assign initialContent_0_44 = 255'h4b29ac56af22e18d40926457dab5aee6f5f9598ea7f0db53bc4e4a94e04f09a8;
  assign initialContent_0_45 = 255'h4d713a79af265adb3877b938b0ae7fd4ad76a6960e8c6f42155106254ed8516c;
  assign initialContent_0_46 = 255'h4e1c057b8dfb64842ba0de58a05289e0b20780457c1a34ec9652b6dbce0d83dd;
  assign initialContent_0_47 = 254'h36f88372c009fc993286d7f40257fc161b060b4a1ca4983b69036e305f87d5bc;
  assign initialContent_0_48 = 255'h50561122dcb9a342cdbc32fb0298da4a6d2923203522169f7b6a3c46293d54ac;
  assign initialContent_0_49 = 255'h73b7860fa6379af73e718277865a3e8d5111532cfb347b625ba5e04b92ad38d7;
  assign initialContent_0_50 = 254'h20056b9fb801dc442db53edcb050696499c7da58d2a653874788912123895022;
  assign initialContent_0_51 = 254'h268ec8894792136915e0adc539329abf24c767ee2295f5df55571a426453b6c5;
  assign initialContent_0_52 = 255'h4e2bd85efc52310851b742c56db7de3ef4cf316a37b54721eb72acc533ecf1a2;
  assign initialContent_0_53 = 255'h4175e26538109ede0800400ba6624b219a042735d6353edae1c7d5464ad1bbd7;
  assign initialContent_0_54 = 254'h23e1291393686042f4dd157fb3c49cdf24c7307f66437989d0ec7a3fb1a49462;
  assign initialContent_1_0 = 255'h4597c2d5e03e62d3de6b94c51cc6e2f7f0363b0e12f1786681f928e3db1913af;
  assign initialContent_1_1 = 255'h5d71428fdf05feb52ab1608cd6f5e16328c4077d48b60874a816abe2988b5914;
  assign initialContent_1_2 = 254'h3862339cef3f4db32ce67758e7377cb7c8d27ef2fc538e7007655c5d6fe32425;
  assign initialContent_1_3 = 252'hb81fb35752a40ad12234eba5807eaecfb79d76992c0e628186bc66979454c85;
  assign initialContent_1_4 = 255'h5d30719d092fa3418884208726c62aca9ae9775ca05941aca20500230a89c43d;
  assign initialContent_1_5 = 255'h4fed9ae55f5cc41e3b53663bf560a30e1f573245dbcc8e60fcd1afe1e4b1a7be;
  assign initialContent_1_6 = 253'h1e5b8b83b9a542b6e410381ff5ce8c263b86b1e9645f63807a1a23a4c10f420b;
  assign initialContent_1_7 = 254'h2ff1c36c1fb11479f5fde194d0ff0330f88c2a9824f96238b7673ec6bc4274e0;
  assign initialContent_1_8 = 253'h16ba36d8d69190005c7d0a7fd56d1296a798cb33fbb7546d9d55ebc6811294da;
  assign initialContent_1_9 = 251'h459fb246e293148529adc6af0e7437222411036404d1738abd6c77b04ed85d7;
  assign initialContent_1_10 = 255'h41b0fb1940ec289c59250f061931bce62b6693bf2781bf67bd65620996c91ac0;
  assign initialContent_1_11 = 255'h5360e84beeb42d5f3c9aa86d70d68392aaaa5879ac7fa63dc4ad7ef4708ed9f2;
  assign initialContent_1_12 = 254'h2afd930d397906bb10c5d03c28ca848e83ae636bada15d5e613298b917a429ec;
  assign initialContent_1_13 = 255'h5874df8d5d1fd55cc73bb91037fb5b9763045c8ebebceec0a222b6acb4563dde;
  assign initialContent_1_14 = 255'h5931eb7da15904697c167ae1b7cd4286399976ffee6a2ea8a71b99e3dc735807;
  assign initialContent_1_15 = 252'hc7dceaff1904c70a941d4d2de10863f8c3a2544be24d6f2119edaea9f361974;
  assign initialContent_1_16 = 254'h263c9da675c9422120f722f46951846ec1f02e9aef10697fdc032cbd56dc83b3;
  assign initialContent_1_17 = 254'h242b82b2e7bf7b9b76ffecb1ff97eea1d3f3678ae85358b5fe94aa89932497ac;
  assign initialContent_1_18 = 255'h64eb9e39284964db76e4e17a787358f089e5e1a2fa6579183237cb0d93c86e22;
  assign initialContent_1_19 = 253'h1d1262ce8246e4bcc1aefa1c6bfca1d0ec43082a46fb3ea78f188b2b206a06a1;
  assign initialContent_1_20 = 255'h4765cccc0995c0b682504648d135107fc1785acccc713c5dbccb53a92ed15f33;
  assign initialContent_1_21 = 251'h466c13d260fd8b9930e655554cc29c2ee7bcf3116902a8429a1d2b461e11b9c;
  assign initialContent_1_22 = 252'hf70d9d2e33b41375d443de27337e5e7c6472a74301e2d9d7963de1b71686d6f;
  assign initialContent_1_23 = 255'h685899a3f56f1a5e5cf0135f77909d7c40ef768d288438b69ca6e00347ada9da;
  assign initialContent_1_24 = 253'h1b7f5e8164db7831fa3ce721522931db555d746891b9a7a4ef88308625da0fe1;
  assign initialContent_1_25 = 255'h5c150bb6c1b1796b49980974d67028230be283db4c6631b6bb132518dc794737;
  assign initialContent_1_26 = 253'h16a801e2ca1bec16b089498c9992d3cb4c7d8bb9a0f8956165ffe9de4ef05eac;
  assign initialContent_1_27 = 251'h440d74e3d73be2a9c2a5721680b983fc52df6c9b486053feb3d3016ec90be2c;
  assign initialContent_1_28 = 255'h506893e963ef99fa7cd8187e4568c91a044fb5287f397151df461353a29ba615;
  assign initialContent_1_29 = 255'h6161a3b78b558aa7c77a19bd48d17a29ac67099939c436a88a1686e33068254b;
  assign initialContent_1_30 = 255'h5781b50088d9b37a391f7f46e6b6174dce8659ac792dc79e205b27abc74be705;
  assign initialContent_1_31 = 253'h1b8bf1984ecf01afd18b0bbf0413ceba2f396c82495b4957503182bc6489d9c5;
  assign initialContent_1_32 = 254'h2a0391b30c3cc24ee2e39a25b4b620d9a5f7941db46b864c992fe097694d4d0a;
  assign initialContent_1_33 = 254'h2dc377e3d7ad99380aca44d812385100fe78ff324ba6d7fc0e67a921303d2f28;
  assign initialContent_1_34 = 255'h6b0971e4d13b1b2ae338c539d9acc17ff46cf9fd2b677b4390ff1a6fc2d66e2e;
  assign initialContent_1_35 = 255'h716a10a5be411170fddffcd38ead5a31da5749b7a87e86573e240f325c9b7b58;
  assign initialContent_1_36 = 251'h775c3d9313c3ebc5f7f952f92fab7b6edc9aa6625498311b2c1fa6a82657ea2;
  assign initialContent_1_37 = 255'h5b6af24ab6887233a3efc2e60691056acf03c93b79ec1804f60e2d293357b0aa;
  assign initialContent_1_38 = 252'h854dc9133532560238a22c7baaa7f1ed55a5aedc5c12dc08c1efe571f35ea34;
  assign initialContent_1_39 = 254'h23d5a01086d25d2575956bee3c94b4a8d064aa6da247cb15f2b3f8bb4cb742c7;
  assign initialContent_1_40 = 254'h2994ae1dcfbb7e488146247f0f7952482a1b84458b14a4e2c88dcd78ef8e8a41;
  assign initialContent_1_41 = 255'h6d46cd37f4f25ca74c96e50bb05f76369feb42b972d577e751b9c6a29d07c17a;
  assign initialContent_1_42 = 254'h3db6370ce200cdb3200475d68b91c405548eca1fe47ef8195c399e3f8dafd570;
  assign initialContent_1_43 = 254'h232a6740632f35ec289f560fb28dc6eeb5b47171bf4a0bde512bbe501beb9633;
  assign initialContent_1_44 = 255'h4394d1b3ca5be52f54d39bb6bc2bda6819cb350346960f7f79c97d7bcd149c7f;
  assign initialContent_1_45 = 254'h2bd3af22c1fdfe91cac8a70bbf722793c3d6e7c253952325d7936bedb1186278;
  assign initialContent_1_46 = 254'h315acb8b0bdbe947f0ceed16b7290dcefdd615eca041fa08327489483312c484;
  assign initialContent_1_47 = 255'h6c4d05497adf2263a2a1bee5e72979d171597c6a7799350a947da2fed08d50f0;
  assign initialContent_1_48 = 253'h10c01c28a57da7a9cadc9c4786d1bf6fb77a76ed693920b9919c890a4a6a077d;
  assign initialContent_1_49 = 252'hbf150f7e34b02ad721a13430fa914fab956cf66adbf94b035f4d040699820f8;
  assign initialContent_1_50 = 255'h6000793141b303a6d7947994fcb43c19487456a795716dece4fda88fcbbfc202;
  assign initialContent_1_51 = 253'h104f6a328d08fd372b3eff88d3cecb804ca4226adde0d8d57bf9157c0d5d38c7;
  assign initialContent_1_52 = 255'h6327fa5e0e5291fac88e8a9f9a4abfdbb2518580227e8094e47a0158baf2b790;
  assign initialContent_1_53 = 255'h56cd2a9097b7a8fcd426bfe372ae3a783ad42da2ddc5abc1f9c8b1a7e777029a;
  assign initialContent_1_54 = 248'he36dd3da1e795fd26da550df4238007d905a43b02659321fa1be93d86e68a4;
  assign initialContent_1_55 = 255'h6b212c40afd2dedc10d055d9c48275aa7ad9a5220a964d48074a093c6375d3bc;
  assign initialContent_2_0 = 255'h719c547de433d29c2aa6ad9d6e80a0fb16f32ef0f3197d50442ed24d7d035b70;
  assign initialContent_2_1 = 255'h5364827a40445fd4cf9d227c5898b763978e94be3b319525893f6a6bb0bd38de;
  assign initialContent_2_2 = 255'h4a64656d98a5d828986a903f37061bd238245a89ebc33130b91bffc36c4e9743;
  assign initialContent_2_3 = 255'h5c91def5f9e7061af94d64da1cba47135262cb105422e7bf1e3964ff5b21f10a;
  assign initialContent_2_4 = 254'h32380af6895cd3c5dc99af8da929f40d5f876296c1ec8bc96c8d608416fd1cdd;
  assign initialContent_2_5 = 255'h54f630a63e7adad91b63c8c5f588c12d4bb232874c7546f5cf447dd7578e38a1;
  assign initialContent_2_6 = 252'h9836e5deed44fe15ff8b65bee710dd4840e211e32eea5edcaa9f55b167d0d90;
  assign initialContent_2_7 = 255'h726652dd154ccfe23dd206f78b2daae991ac284007c172f4d4b89b9b1adb4098;
  assign initialContent_2_8 = 255'h7343f3b646888d89671fe764a77b6799b99359307ee583be10b4bf4c1646bab0;
  assign initialContent_2_9 = 250'h3c992dfe1c2cb83856467ebf83426286b7ae65e6336ae3c91ff1d398ae0de67;
  assign initialContent_2_10 = 253'h1c0eb0a1eb09022e5882d04f17b58d665fcca167bf926683eb8b0200d51d1d61;
  assign initialContent_2_11 = 255'h5b78b552b150025bf4dc5f74f7187bb95f1c625216408aac36b25f93aac824ad;
  assign initialContent_2_12 = 255'h409d072638627609c116075527e3021e35e2f7a45a72c89ccfdb0f3ce8ac1dd0;
  assign initialContent_2_13 = 252'hf58b72cdef8c4f7da9b732e6e67fe6991e3b248e5114b8d7c3a48b87215230d;
  assign initialContent_2_14 = 253'h18d6ed4cb9bd646d0f01fdaa90e044ad44122c4d33cdca2f355397a386deda10;
  assign initialContent_2_15 = 254'h28327d51f6723b41923a154f3647362ce549ace26c29ba658dc00c22c7265e5a;
  assign initialContent_2_16 = 254'h278d6a97675fd062938bd33df3c17f2eac780af52e14e068c7f906adc777da1c;
  assign initialContent_2_17 = 255'h6853c380081f1de555ddd016eb9449723578397bc342a5a1ab50deeff2e6666f;
  assign initialContent_2_18 = 255'h43901fad86a42bbdfc03a5380496b1ae2dbcc848218c9df3e9a89c86ffcfd706;
  assign initialContent_2_19 = 254'h2fdf2d02ba2614843da21bc7d15751e1e14c7e8939f060e8a77544898a964787;
  assign initialContent_2_20 = 255'h4919468964d0adfe78b0b03874005c682514a271964005477ffe51cddae33fe1;
  assign initialContent_2_21 = 252'hbed0481c1d3a1cfa93a234548d236f07eb9974f4fc118a427a4906e15bff10b;
  assign initialContent_2_22 = 252'hb1f43ebce8274c63b498e9afb08d7db5d6c461dec6ef7c430bd8a70325e1a5b;
  assign initialContent_2_23 = 253'h166bc3586286bc195d562323ccb3f2767464fd4adf17b145428d56d1a3ebcdbd;
  assign initialContent_2_24 = 255'h682c01c08691ca5398e21766de998908d97cd2693488b2dc77dd98fa93ded68d;
  assign initialContent_2_25 = 255'h55e3675cbde7b7f54a8542889e7e08c69b73f929833e99d2f8eafec229aef400;
  assign initialContent_2_26 = 255'h6c0cf0f6608d9dec58faaa544dae05cb9e4e8b551757e37b060be016f4e04f28;
  assign initialContent_2_27 = 255'h44db06be530ddf5fd0c7617d941532b0e18760fc527c80bb7b35c8bcba79f102;
  assign initialContent_2_28 = 255'h64228dc41a1daa01d70310233b00fe449382f29f034efe1dd1d270b8dd5d4e2c;
  assign initialContent_2_29 = 254'h3e23f72361d9564ee642fa245bacd1ad5c2fec3353bda0126d39eb87848b7693;
  assign initialContent_2_30 = 255'h5113fbb31d3a7b50ad7563dfd9180253982d04b77ba0d270368de730f1c2d142;
  assign initialContent_2_31 = 254'h2ca9282e5e798ccc5c46aa9a27c5c63d1c82adcec28afa87c2def9debbfb0423;
  assign initialContent_2_32 = 252'he816050f009975e9b5c5a761b66f6897952690276fd05815dadbe91113b3f2f;
  assign initialContent_2_33 = 255'h40e1ed7492a10495b5f3443153887f2f1e920196016bd50415fe657fbd445090;
  assign initialContent_2_34 = 251'h4ec0186bf9baba76703ea27f4fc06ad1c08b181bc62a49ca0b7bbf151df66de;
  assign initialContent_2_35 = 254'h23c5d71ec7f1f19638fce402907c5643e29cb5098f0fa87b58850675fb6d7bd8;
  assign initialContent_2_36 = 255'h50f7d37aeee78a630aecc3cc5017a812943e903205209696107599496e3bff23;
  assign initialContent_2_37 = 254'h21e421bc6c570eb53a56a45c4ada293fefe3ed0f115263bf502981cf8d6a64fd;
  assign initialContent_2_38 = 254'h368ae1626461f6d9a5a35888060d38e61498d047da74b55f3134f65363989975;
  assign initialContent_2_39 = 255'h412c09ebef9a00dde8facc0fdcc2f89fec4a877001a22d35cabf975136c304de;
  assign initialContent_2_40 = 253'h1cf89973996e33a5432b15595ee19cf2f50ba4facc15b5a49162285784517a31;
  assign initialContent_2_41 = 253'h1be13383c54535d3431242bc2d4cee22b109d9d8d80df846b891604de2a69f0f;
  assign initialContent_2_42 = 254'h275c1332218c4221e3cd1382f4580c3740c4d64fc475e51dd533eb828c711955;
  assign initialContent_2_43 = 255'h44cbb1b0e2d216081aa33593d10ea35a89091e201cef6b243dffe9a3a9cc6d2a;
  assign initialContent_2_44 = 255'h6d87561e194eb0aa03d8c86b2b3638ea099216e25dac662209ea098177a1f012;
  assign initialContent_2_45 = 255'h5548a2cb6494202dc9ccd53c28a646e380f33a77bb27acdd409a2a608c0bcf31;
  assign initialContent_2_46 = 252'hafd0c8d17c218fa0f606909a6f6b9ae50b097acbfa9e3ad981b87b7df5d50cc;
  assign initialContent_2_47 = 255'h57222e019a99df6e8b86c1b64388ce068d0e01d9cce358f678da35dfe86639a1;
  assign initialContent_2_48 = 254'h3f8bec0774d7dd76f945e363e04bac528631708c620c374821924216112283cc;
  assign initialContent_2_49 = 255'h4aa90213015df3c5a3de82935129270a95c3cc0abf37d81501e98db745d7cf27;
  assign initialContent_2_50 = 254'h3839dfcfc80a2d9c3ffd971c75c52ff2fda7ce7b03b7d105d9ca5ffdec654241;
  assign initialContent_2_51 = 252'hf2b3adfb545911a3f459506fb4cd03607d6082726e8fe24e521e3836f02f4b1;
  assign initialContent_2_52 = 254'h2d9efdd3811a9cb5d04c7e2fca02988e5021d03fa91bb6ded940caae7955e54b;
  assign initialContent_2_53 = 255'h5f259c25fb57b0cb9f13c32e3c5010d6d36d69c14dfe7f9fbeb04b1d9504884f;
  assign initialContent_2_54 = 255'h5acafa8f5c9e614f236eb89ea6682ffd819bbe5cc61430dc5140afbcb91cf4ad;
  assign initialContent_2_55 = 254'h3d12c6e84485a1f8019ffa5efacc5f2bf90b775697c443b8396f6c2862b13941;
  assign initialContent_2_56 = 255'h581f16e55cdfa35319dd21a68aeb6c0ea3b2423e6dfbdfda00e331dad3285027;
  assign initialContent_3_0 = 255'h61ddbd21aa3cdf60f8db05bdee3a2270738e9b1f8233d80246ab0d8ff64b9ae6;
  assign initialContent_3_1 = 254'h3d28bbbe6a5d5f27d1036aa42a4f08bee0107d3d714d9c299419bbbd33e913db;
  assign initialContent_3_2 = 254'h39899330c9a40e0b903eaa430bf4941e82ee5aa3a0ea91f07952fcce3bd19d34;
  assign initialContent_3_3 = 254'h366b123e3d009276b1d843f4e7c56bc8868326c2d705ab0dc7fa011f0beaa92f;
  assign initialContent_3_4 = 254'h3bc0dfe7e55ddb0d5c59e4e91394e9ed01ea7126a450fbdc5ed09de7e3999523;
  assign initialContent_3_5 = 253'h1a01537b2edec1b6866842e5aca0fd6036611a188c4b234bb25a66589d1aacd9;
  assign initialContent_3_6 = 255'h5bdbedf19519efc31383e5b7bdc2b2e43a8c9319943132f71c0704b5f20b5333;
  assign initialContent_3_7 = 255'h49c4a7264eff8c8a35b5566a432f3c878aea939774d5331beb19873433ff5958;
  assign initialContent_3_8 = 255'h6e76c43ce3e34074519ecc717f44cfa4b9904d9336af969d622f45ef3b6c7ea8;
  assign initialContent_3_9 = 255'h6c089cf205db963adeda7f87439955a53cfa2e1d04ca2a76f175565217e90264;
  assign initialContent_3_10 = 255'h53dcab90596ec843142185dda9bca22d9560df65d6d25cceb7fc30347c8f5c73;
  assign initialContent_3_11 = 250'h37ec57a1b4a47f75f2116dd47b888c13542168dc9ebdf3a4f328b9bcb287e4d;
  assign initialContent_3_12 = 253'h1186f410ffdfa0d4976ebc0a580107be377ab9ecc210a85d9881c3f64974d0a6;
  assign initialContent_3_13 = 255'h5d07a354e5ca8788127994b6201c9a2456b5bbbcd04f1fc37dfeee072a67d887;
  assign initialContent_3_14 = 252'hf68a6d19696c4d1c9f0b4149dab96b18e061f651ba3f30554d31f32671ac438;
  assign initialContent_3_15 = 249'h1f8a70d0a5ac286cdbe0f4df7cd134ac27d17873dcfad2753c9087852b396e4;
  assign initialContent_3_16 = 255'h6dab0c6c36dabb98b0d0843e25023ab59469dd99d413f13d19286a7126394e97;
  assign initialContent_3_17 = 254'h3426f66a0ded8fbeaa176c5720b13e79c06a8520ad9c4f144c2e39e82f2a3776;
  assign initialContent_3_18 = 254'h2a5002dd7dd294a70c840e4ac359acf9ca296f0c3c5ba1b65077e17b955b9205;
  assign initialContent_3_19 = 253'h1897c311109acfc300dbb0eeccb7c4c571d84e8c989161a3ed94442deb1fcbd7;
  assign initialContent_3_20 = 252'hbee4ca4bfa1aa02c474d7ae19ea04f5b89aaa7f42c184ea96f2131d35afa360;
  assign initialContent_3_21 = 255'h4fc8c2b7c94170a43056b066c48c70a15da307c534f8bcefcbc9a8e8ce7adce4;
  assign initialContent_3_22 = 255'h69878703e3ad4df912cae7ebbb8e04a7d37a8cf90ad4a7fbc05019aebea7f4b7;
  assign initialContent_3_23 = 255'h50650c96e3514d7bca9b9ca6d0ef92de44bd3e564edae4c2da2caabac6f930aa;
  assign initialContent_3_24 = 254'h343e7206996630a936aed8295150695c9fa21e2ae48e2489e350bed59aeed90a;
  assign initialContent_3_25 = 255'h71fd75fe89872cdb69151a1f5d26537e6105162c0dd84abf75136495cf25912b;
  assign initialContent_3_26 = 255'h41fd9f218d0061418d17b1762d562465284070d8add6e161f0e54549d4981d35;
  assign initialContent_3_27 = 255'h5afef959754485e1953640ef55945748e2539aa33a368aad26ffd9786af9394c;
  assign initialContent_3_28 = 254'h2c1a2004be2e92bb3a334ab7479fdf77aeae26aad699d6d3cf767eaeecc91fd9;
  assign initialContent_3_29 = 255'h5732893412d50959c8f56d731f00bbf313c18c693f87f3a513ef9311faaf5c96;
  assign initialContent_3_30 = 254'h337de782119e1928eb44f40de52c719c9723d939d4e0c91dc74cf253b3b2b9eb;
  assign initialContent_3_31 = 255'h4cd303643ea2530f2fc0f00a660654daaad9386bca098e75759fd121eb003922;
  assign initialContent_3_32 = 254'h21e75a288129097d11568099d4d75bcbbca53a1e2c8fe8ad6121b82deed4475e;
  assign initialContent_3_33 = 254'h350580ff40b1a560057c876f70cbb5b4cee6169429af76ba32b201ed9034ff41;
  assign initialContent_3_34 = 255'h5ba3bfca86781caea27395021aff7619922741afeadd381908382dc1cf3a201b;
  assign initialContent_3_35 = 254'h224f10dc5a9e59329be2fe0e57ba3dba53e8148fb143511b8e45e18553dcff80;
  assign initialContent_3_36 = 253'h108f95df62fc095442bc17c8eefd2dab965c85e314309b212d7dfe1aa7d58f47;
  assign initialContent_3_37 = 255'h44ef434d0ee752fc6eb1e3ee1d35415272b8547fda5d1b11ec816b8d179e8f23;
  assign initialContent_3_38 = 255'h5ecbce3cfa879f1e3463ae780f577aa6f7ef8406777af2af4fc83ba504d3fa91;
  assign initialContent_3_39 = 255'h6181c724431ea1591283191d96d0bfc409f008def9ee5dac77e362d27d50dc96;
  assign initialContent_3_40 = 255'h6cdee21312112696fb9815b2af5196a578424707e3fd622449ef24c8e269b1d3;
  assign initialContent_3_41 = 254'h33f75fbee6faaec4c017e01666e82c41d14caf3c13eb047cea2afa40f65cacd5;
  assign initialContent_3_42 = 255'h6f7e6ac9be53cc01f4a27c47418029d2356f0f0b1dd49a231577594af1cd914d;
  assign initialContent_3_43 = 253'h1637226aee56fcb110a7c56a5c08d94a1e509483900129d7af581cb99fb690ad;
  assign initialContent_3_44 = 255'h52c17e35ef264a191039b4adcda8b6ae71127d135428906cc0cadceae2010e24;
  assign initialContent_3_45 = 253'h1951f367c0d8425fbf2e1223608a9647725919f5423a0256f0cfc274f94c2b22;
  assign initialContent_3_46 = 254'h21c39ab35355280b42d7c04613362cb2e8e174cd04e442c05158106cb86d5372;
  assign initialContent_3_47 = 250'h2a72d3b6a083d157ea501dc797f5a2eb3353845aa722dc4c5c251cef0186550;
  assign initialContent_3_48 = 255'h6e45cbb08375c1377dc4fcde17aa183f7fb33851ba6b660b07d7aee44934415c;
  assign initialContent_3_49 = 254'h21f57fbe766addd5fbcb66e39b3ba311da4b03a35219030033a9b419f8445b96;
  assign initialContent_3_50 = 254'h2318c472d8c802c15d668d800f43cfc479a6830c6b2d82c7732ca497f209a11e;
  assign initialContent_3_51 = 255'h596972f4da5a229801a42837661ab63c0485bef98312a90570df72d902190584;
  assign initialContent_3_52 = 250'h2b4bc4cfc6e1b9d4910482c0de050cf42806d3b9d83940e8d93f0b27abb2c1a;
  assign initialContent_3_53 = 254'h2a9a3184aa49ba84200bfff22bce8bd0336eaba598c61fc5e050565e6718f390;
  assign initialContent_3_54 = 255'h64d8caebd3302ee45d49f2a7dbdc40c5d70105649d6714216d862ccf90ff5e4a;
  assign initialContent_3_55 = 253'h1cbdf93c411d6a4aea04b0fc1eb2b1c7b0aa3cf0335430a34614fbff8a5bd71b;
  assign initialContent_3_56 = 252'hf6bf8b42ad4f9f22cd37279f26c5f8852f650a34dda16facea181c8db9bd59d;
  assign _zz_memOutputs_0 = io_partialRound;
  assign memOutputs_0 = _zz_constantsMem_0_port0;
  assign _zz_memOutputs_1 = io_partialRound;
  assign memOutputs_1 = _zz_constantsMem_1_port0;
  assign _zz_memOutputs_2 = io_partialRound;
  assign memOutputs_2 = _zz_constantsMem_2_port0;
  assign _zz_memOutputs_3 = io_partialRound;
  assign memOutputs_3 = _zz_constantsMem_3_port0;
  assign select_0 = (io_stateSize == 4'b0011);
  assign select_1 = (io_stateSize == 4'b0101);
  assign select_2 = (io_stateSize == 4'b1001);
  assign select_3 = (io_stateSize == 4'b1100);
  assign _zz_io_constant = (select_1 || select_3);
  assign _zz_io_constant_1 = (select_2 || select_3);
  assign io_constant = _zz_io_constant_2;

endmodule

module FullRoundConstantMem_3 (
  input      [3:0]    io_stateIndex,
  input      [2:0]    io_fullRound,
  output     [254:0]  io_constant
);

  wire       [254:0]  _zz_memInst_0_port0;
  wire       [254:0]  _zz_memInst_1_port0;
  wire       [254:0]  _zz_memInst_2_port0;
  wire       [254:0]  _zz_memInst_3_port0;
  wire       [254:0]  _zz_memInst_4_port0;
  wire       [254:0]  _zz_memInst_5_port0;
  wire       [254:0]  _zz_memInst_6_port0;
  wire       [254:0]  _zz_memInst_7_port0;
  wire       [254:0]  _zz_memInst_8_port0;
  wire       [254:0]  _zz_memInst_9_port0;
  wire       [254:0]  _zz_memInst_10_port0;
  wire       [254:0]  _zz_memInst_11_port0;
  reg        [254:0]  _zz_io_constant;
  wire       [254:0]  constantsMat_0_0;
  wire       [254:0]  constantsMat_0_1;
  wire       [253:0]  constantsMat_0_2;
  wire       [253:0]  constantsMat_0_3;
  wire       [251:0]  constantsMat_0_4;
  wire       [250:0]  constantsMat_0_5;
  wire       [251:0]  constantsMat_0_6;
  wire       [254:0]  constantsMat_0_7;
  wire       [254:0]  constantsMat_0_8;
  wire       [253:0]  constantsMat_0_9;
  wire       [254:0]  constantsMat_0_10;
  wire       [250:0]  constantsMat_0_11;
  wire       [254:0]  constantsMat_1_0;
  wire       [254:0]  constantsMat_1_1;
  wire       [254:0]  constantsMat_1_2;
  wire       [254:0]  constantsMat_1_3;
  wire       [253:0]  constantsMat_1_4;
  wire       [254:0]  constantsMat_1_5;
  wire       [251:0]  constantsMat_1_6;
  wire       [254:0]  constantsMat_1_7;
  wire       [253:0]  constantsMat_1_8;
  wire       [254:0]  constantsMat_1_9;
  wire       [253:0]  constantsMat_1_10;
  wire       [254:0]  constantsMat_1_11;
  wire       [251:0]  constantsMat_2_0;
  wire       [254:0]  constantsMat_2_1;
  wire       [254:0]  constantsMat_2_2;
  wire       [254:0]  constantsMat_2_3;
  wire       [253:0]  constantsMat_2_4;
  wire       [252:0]  constantsMat_2_5;
  wire       [254:0]  constantsMat_2_6;
  wire       [253:0]  constantsMat_2_7;
  wire       [253:0]  constantsMat_2_8;
  wire       [248:0]  constantsMat_2_9;
  wire       [253:0]  constantsMat_2_10;
  wire       [254:0]  constantsMat_2_11;
  wire       [254:0]  constantsMat_3_0;
  wire       [252:0]  constantsMat_3_1;
  wire       [251:0]  constantsMat_3_2;
  wire       [253:0]  constantsMat_3_3;
  wire       [254:0]  constantsMat_3_4;
  wire       [254:0]  constantsMat_3_5;
  wire       [254:0]  constantsMat_3_6;
  wire       [253:0]  constantsMat_3_7;
  wire       [254:0]  constantsMat_3_8;
  wire       [250:0]  constantsMat_3_9;
  wire       [253:0]  constantsMat_3_10;
  wire       [252:0]  constantsMat_3_11;
  wire       [254:0]  constantsMat_4_0;
  wire       [254:0]  constantsMat_4_1;
  wire       [253:0]  constantsMat_4_2;
  wire       [254:0]  constantsMat_4_3;
  wire       [254:0]  constantsMat_4_4;
  wire       [254:0]  constantsMat_4_5;
  wire       [254:0]  constantsMat_4_6;
  wire       [254:0]  constantsMat_4_7;
  wire       [253:0]  constantsMat_4_8;
  wire       [253:0]  constantsMat_4_9;
  wire       [249:0]  constantsMat_4_10;
  wire       [253:0]  constantsMat_4_11;
  wire       [254:0]  constantsMat_5_0;
  wire       [253:0]  constantsMat_5_1;
  wire       [253:0]  constantsMat_5_2;
  wire       [252:0]  constantsMat_5_3;
  wire       [253:0]  constantsMat_5_4;
  wire       [254:0]  constantsMat_5_5;
  wire       [254:0]  constantsMat_5_6;
  wire       [254:0]  constantsMat_5_7;
  wire       [253:0]  constantsMat_5_8;
  wire       [254:0]  constantsMat_5_9;
  wire       [254:0]  constantsMat_5_10;
  wire       [252:0]  constantsMat_5_11;
  wire       [254:0]  constantsMat_6_0;
  wire       [252:0]  constantsMat_6_1;
  wire       [253:0]  constantsMat_6_2;
  wire       [254:0]  constantsMat_6_3;
  wire       [253:0]  constantsMat_6_4;
  wire       [254:0]  constantsMat_6_5;
  wire       [254:0]  constantsMat_6_6;
  wire       [254:0]  constantsMat_6_7;
  wire       [251:0]  constantsMat_6_8;
  wire       [252:0]  constantsMat_6_9;
  wire       [249:0]  constantsMat_6_10;
  wire       [254:0]  constantsMat_6_11;
  wire       [2:0]    _zz_memOutput_0;
  wire       [254:0]  memOutput_0;
  wire       [2:0]    _zz_memOutput_1;
  wire       [254:0]  memOutput_1;
  wire       [2:0]    _zz_memOutput_2;
  wire       [254:0]  memOutput_2;
  wire       [2:0]    _zz_memOutput_3;
  wire       [254:0]  memOutput_3;
  wire       [2:0]    _zz_memOutput_4;
  wire       [254:0]  memOutput_4;
  wire       [2:0]    _zz_memOutput_5;
  wire       [254:0]  memOutput_5;
  wire       [2:0]    _zz_memOutput_6;
  wire       [254:0]  memOutput_6;
  wire       [2:0]    _zz_memOutput_7;
  wire       [254:0]  memOutput_7;
  wire       [2:0]    _zz_memOutput_8;
  wire       [254:0]  memOutput_8;
  wire       [2:0]    _zz_memOutput_9;
  wire       [254:0]  memOutput_9;
  wire       [2:0]    _zz_memOutput_10;
  wire       [254:0]  memOutput_10;
  wire       [2:0]    _zz_memOutput_11;
  wire       [254:0]  memOutput_11;
  (* ram_style = "distributed" *) reg [254:0] memInst_0 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_1 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_2 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_3 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_4 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_5 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_6 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_7 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_8 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_9 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_10 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_11 [0:7];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_0.bin",memInst_0);
  end
  assign _zz_memInst_0_port0 = memInst_0[_zz_memOutput_0];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_1.bin",memInst_1);
  end
  assign _zz_memInst_1_port0 = memInst_1[_zz_memOutput_1];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_2.bin",memInst_2);
  end
  assign _zz_memInst_2_port0 = memInst_2[_zz_memOutput_2];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_3.bin",memInst_3);
  end
  assign _zz_memInst_3_port0 = memInst_3[_zz_memOutput_3];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_4.bin",memInst_4);
  end
  assign _zz_memInst_4_port0 = memInst_4[_zz_memOutput_4];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_5.bin",memInst_5);
  end
  assign _zz_memInst_5_port0 = memInst_5[_zz_memOutput_5];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_6.bin",memInst_6);
  end
  assign _zz_memInst_6_port0 = memInst_6[_zz_memOutput_6];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_7.bin",memInst_7);
  end
  assign _zz_memInst_7_port0 = memInst_7[_zz_memOutput_7];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_8.bin",memInst_8);
  end
  assign _zz_memInst_8_port0 = memInst_8[_zz_memOutput_8];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_9.bin",memInst_9);
  end
  assign _zz_memInst_9_port0 = memInst_9[_zz_memOutput_9];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_10.bin",memInst_10);
  end
  assign _zz_memInst_10_port0 = memInst_10[_zz_memOutput_10];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_7_memInst_11.bin",memInst_11);
  end
  assign _zz_memInst_11_port0 = memInst_11[_zz_memOutput_11];
  always @(*) begin
    case(io_stateIndex)
      4'b0000 : _zz_io_constant = memOutput_0;
      4'b0001 : _zz_io_constant = memOutput_1;
      4'b0010 : _zz_io_constant = memOutput_2;
      4'b0011 : _zz_io_constant = memOutput_3;
      4'b0100 : _zz_io_constant = memOutput_4;
      4'b0101 : _zz_io_constant = memOutput_5;
      4'b0110 : _zz_io_constant = memOutput_6;
      4'b0111 : _zz_io_constant = memOutput_7;
      4'b1000 : _zz_io_constant = memOutput_8;
      4'b1001 : _zz_io_constant = memOutput_9;
      4'b1010 : _zz_io_constant = memOutput_10;
      default : _zz_io_constant = memOutput_11;
    endcase
  end

  assign constantsMat_0_0 = 255'h489ac9289b121784c79133e51917e24610abda74708f0f48656e5817de651e01;
  assign constantsMat_0_1 = 255'h6aae617b93294ecdcfcf0e578c5681dc7ad383cdbace5474d6269493b756e4f8;
  assign constantsMat_0_2 = 254'h259af037a7e7c5fde581f4601d23f681dfc1a92f028cdb1318ebdfd7fcfc2573;
  assign constantsMat_0_3 = 254'h26b8e174187543023c9f463f2b4759028c3d3090380ad7da7f3b5f13c8238b86;
  assign constantsMat_0_4 = 252'hc2b6b23e1d9f4c34f338e85bef39f560a771d31d8e8f911dc5b589415204a35;
  assign constantsMat_0_5 = 251'h4f7f4eebae9aa0f4d6ac4b0111efbbf61bde34e854741ff9431dda4c402733b;
  assign constantsMat_0_6 = 252'he5e22194181e51c9f22478d53e43776fc65924743eaaab12b1f4957cb8d87c3;
  assign constantsMat_0_7 = 255'h5ad01fd9949dd1951e53cb7df7be004c344fd0a1685497edc8dbaa61a4e0157e;
  assign constantsMat_0_8 = 255'h66b3e16e1da5ac4e9d70e35e54fa6f268883334f116147b79574d0f05065820f;
  assign constantsMat_0_9 = 254'h2709e8dfaa6acabd0c665fddbe7f467d7bfca5100fef26a0015a32963414a372;
  assign constantsMat_0_10 = 255'h67d4d856c7c8a939022ea6ab3061e1f5e103092bcb73d637c030821561a48dda;
  assign constantsMat_0_11 = 251'h7dcb5d1869b0ea4e804cf5aef01787c79ccedfc91475f0d804bfc487490e42e;
  assign constantsMat_1_0 = 255'h47f04a041bdafefa028db1fe28e08b6a13cea63cc0b9d3f2320842475bdc8ae2;
  assign constantsMat_1_1 = 255'h737781762f6972ea516174a0d45fc0e6e07d7bd2674b59b45136c27eb21506df;
  assign constantsMat_1_2 = 255'h638221e89540eccebc26f3ab0b2e91180db55f2665cb7bbbf9ef761623009b7e;
  assign constantsMat_1_3 = 255'h4b74b782be2a6336ff8d7f37b2ac091bb35e77e53e5cc798c95191fdae2f5a86;
  assign constantsMat_1_4 = 254'h325dc076a94d627905cfa6a771e73262a7e465a69bbac84f19e75078dbc66f90;
  assign constantsMat_1_5 = 255'h53bc3c14c92c6f98f9d726617e805b6d8dd46a0ca65623fe2a95f91b06ac71fe;
  assign constantsMat_1_6 = 252'hefb5f9c645afe1975067561958d6e2dfe51a49209ca1b18478f73aac4a7edf4;
  assign constantsMat_1_7 = 255'h6f8032f43ab561f86c796cf6242e53283e433c373d91a9a35f5b138c297d0f61;
  assign constantsMat_1_8 = 254'h2c2f07fd44b8e6996b0af65d7e98d8bd95003f11635160386d2331f882254573;
  assign constantsMat_1_9 = 255'h488d8a4f3ecbcf6b47874cf1cc18eb6965aeca29dc87f74e607138f005e23d25;
  assign constantsMat_1_10 = 254'h3b82233053b0f782eb5d94560c60edf554f26b623fc50a2111f94ff2e08d88cb;
  assign constantsMat_1_11 = 255'h6cb359e9802cc97add5749bcb82cff9d480725fbcee27d040b11ee53282d557e;
  assign constantsMat_2_0 = 252'he048cb4a14e76c48aa7c94bcb62eefab1d6cd81535bc6da2fae43c9d5dce3c0;
  assign constantsMat_2_1 = 255'h450c8bdfdb1b3bb48c42c03de7156f5463d145ebb724e5cc46407b8cc0274e50;
  assign constantsMat_2_2 = 255'h52466d9dd56dd54d40c4243c2aa7c1b973ca36d9a861dd456481bd1cb2e62b84;
  assign constantsMat_2_3 = 255'h49346ac358b17211f95da95826b3af84c91586eb6a6b1ca93c4667bec8d58587;
  assign constantsMat_2_4 = 254'h3109c0e791242e656446a280f2f3d45d44a7f2faada7633af8bf16c5663d3917;
  assign constantsMat_2_5 = 253'h13b40fcacd8a5f5b661604a746dc189193f04ac0346fa9c40ba94c2699051d78;
  assign constantsMat_2_6 = 255'h606db33ea58b35ad8cc4e5a5227d7cdbda1d519c79ce33e240e645ff350c144d;
  assign constantsMat_2_7 = 254'h2eac2753a1b1db26b2e0e12569cb113af2e6315dffa1711d2577505ff577c88c;
  assign constantsMat_2_8 = 254'h2c2dd0296cb307c11b987bcd415515459480a1c77111275356e9f6e631d19d17;
  assign constantsMat_2_9 = 249'h1a19de7191292d6e57df4cf46ef2a7db4215c4bde7e3769dfcddfd749a67690;
  assign constantsMat_2_10 = 254'h384dafd721307dd80af448f34cdfb1b81e43adee3b245a96329bd2bc47dc34c8;
  assign constantsMat_2_11 = 255'h64c241c5f35e4c954545e0cd58f265e5cca991a186c11c9392d87e06ffd24b81;
  assign constantsMat_3_0 = 255'h673805124a7f8e5d015e25bfdb0a4c683ca5edd130fb9bd31910eb5e2c06b121;
  assign constantsMat_3_1 = 253'h1ac35e27f873308601736fed0bf0905ccc323a2a4806ddf5053eb0e3165d2241;
  assign constantsMat_3_2 = 252'ha10fd5975766908c77d390b886e67a10a5ba942d7aa6a2728b7dba89c631d2d;
  assign constantsMat_3_3 = 254'h202a4693c0984afc439478399a0f8d41d836c4c253305b074bad18b6636215ab;
  assign constantsMat_3_4 = 255'h407ccd54e212084ec86c455c47abf8ea44fa2058257cb6da6795bad57334af59;
  assign constantsMat_3_5 = 255'h55943894574d996c9a599f6c0cdc040b63c9474d7f11b326a86ae5c4a56334b2;
  assign constantsMat_3_6 = 255'h40dfa76f81e1bd61266dfc8d56c436bf4e8ce6619d5bbb983e29a36bb0ae04a0;
  assign constantsMat_3_7 = 254'h2f8f3d8c07d30b2a5ccb8c330804836af8e600420c4802b9296af604b4cef7f6;
  assign constantsMat_3_8 = 255'h55ee7303d0121e0c4475da2ddbffb0f389f250e431829c2dad74a6b9b2ee4e13;
  assign constantsMat_3_9 = 251'h655178cd78ba47238f713c590ec999a3395e0045828d6686601b47d6f8eb2e6;
  assign constantsMat_3_10 = 254'h3b01c21370e105db41e5affe4786633f6c00b9a5e6295f0bad0db63805b0ca9a;
  assign constantsMat_3_11 = 253'h13e01879b679f68fcbff6dbe7c8923a4a1ea5fa4e8ccc9a218502b8d12255df3;
  assign constantsMat_4_0 = 255'h4d4496eb98eab7e3e1bbb45428f95c5d400026f4bfdb95013c747146ae977273;
  assign constantsMat_4_1 = 255'h701099c099cfde2096e1f869921804a6c70b4ac4274ee5c7e35c6aaa696400b2;
  assign constantsMat_4_2 = 254'h38954be1c280b0711ff40645893b7be84a4181382c0dc9551dfca9fd466305b9;
  assign constantsMat_4_3 = 255'h53ab2b1c5875ec882702051a1a8f1be98fe5bbad2ba3f88ee83a653c9399a482;
  assign constantsMat_4_4 = 255'h5e9a34ad9154a78f6f5aa86e4675c881aa2e7f369c0c0512cb2656ad306f8523;
  assign constantsMat_4_5 = 255'h435d51dc5b123ac7604f07fefba091579ccd4f8d5de048f31dc0ae4c117ac9ba;
  assign constantsMat_4_6 = 255'h65bb6803d56f0643476becf7885f0838439db8ea4b142298028548e0195a751d;
  assign constantsMat_4_7 = 255'h4500a30faf31f2bba4a34da9d27ee679b756a441704ee0bc51ebd349b0898034;
  assign constantsMat_4_8 = 254'h39c0ec5521a70d19d15bcef222e5289ed2f9b8a86b3df23639202b951264b2d8;
  assign constantsMat_4_9 = 254'h26d48fa2037d87d7287acd9decb6cc182ccd14151fe2e4aa39e122635d38d1a0;
  assign constantsMat_4_10 = 250'h2f485ddfe7dcf99bc738c8dd2833d02e713c7996b4ece52d69574d5f2e4ce42;
  assign constantsMat_4_11 = 254'h34deb0897d57fd35e7640d7d0ef34b33d0d65e72d8e242b78bd80181a5badc73;
  assign constantsMat_5_0 = 255'h45ceb97c8e0e7586c3a7393cadb7ddfaa33c05cf81307364f41e541d41f1cb0f;
  assign constantsMat_5_1 = 254'h3f44295c4a1438722922df6acebd4168802b977626d942653b741423ba9b69af;
  assign constantsMat_5_2 = 254'h2eae724b7c053bb8250cda3b57a79293a3d707a37c0a66a07ca178f29fbf803d;
  assign constantsMat_5_3 = 253'h1e64207bbd21cf35b632ca8c90fb340da4067fa165849580b495009fd575bc36;
  assign constantsMat_5_4 = 254'h3e5fcdfc0b606afe6960ad5b8afd1e7baaa47cb5b6bbfcdb71a442e7985776ae;
  assign constantsMat_5_5 = 255'h73978eb19d784b11350e95d51bf198337d723ea813248769ba99322a31363da0;
  assign constantsMat_5_6 = 255'h6ecb03831f4d1c30d9aa59db5b13664a741fcb551e49dfa6e45d5b11af6d1f84;
  assign constantsMat_5_7 = 255'h56417a4978f1949eab9685ec80c94a9b751e8254d74013fcc2d4757128537005;
  assign constantsMat_5_8 = 254'h3abc30c9d794d437f34d8d4ab470398330cbfda0a67018e51df762deea9d3068;
  assign constantsMat_5_9 = 255'h5b78e2c3427b3499b1f636fb275491f767ee60ba238c185c8bd1eaa6692eb84f;
  assign constantsMat_5_10 = 255'h736543df297e26944470d01bdce64b17f8a11d50ddaf11243628e7fa0e1614e9;
  assign constantsMat_5_11 = 253'h144b278b192092f241f894c055b157d491be170beea68d3647fe8f3cb945279c;
  assign constantsMat_6_0 = 255'h6e5a17aabb6838f38171fbd2675c1eed7c7afb1c046e65860401819a3374b0f8;
  assign constantsMat_6_1 = 253'h1d4b037dec167f9b9e98018fe50c9fe7627ee72a90d7c995b1784bc99713871c;
  assign constantsMat_6_2 = 254'h317de90bd5946fb28e525ede21248a0a9203fcef8cf15eec45cba75ca4541558;
  assign constantsMat_6_3 = 255'h6fab7fb4718b40810ebf39b39a01ac641cb57c455829949d59dcfe51745c1560;
  assign constantsMat_6_4 = 254'h2da3c9986f6250ca25d6ce3e2053c81ac7937d924acd31f1c3915b4bb678e8bc;
  assign constantsMat_6_5 = 255'h64d69fc29cf0bfe8ec8ebf22e46575df5505c78799a637d1eb5f25ec1f3a582e;
  assign constantsMat_6_6 = 255'h4a8cca333a0d60a5d014f5f3fdfe73f4c9f55a1674e897ddb1a416bfa22cf2df;
  assign constantsMat_6_7 = 255'h5f2eaa1e0658efa57b0f2096f590d9d7b32b0c9dc797590cc89e820f8f88023b;
  assign constantsMat_6_8 = 252'he0b21be246a9cb838939c8f3faaa96afdcb571a274305dda5ccdf8b6109894e;
  assign constantsMat_6_9 = 253'h1d84b55d20c7e0c7c4cf89b3102bfa22a07f62362d3fb125dd0c1a2f12888521;
  assign constantsMat_6_10 = 250'h3f3d0f2a6ec1698e1df3931e9d487caeb58a4f04065fe5f714964ba04df671e;
  assign constantsMat_6_11 = 255'h625c6847a00daf49fee2b25a8494ad6ae045940c2c33ecf17284a942f1198bd3;
  assign _zz_memOutput_0 = io_fullRound;
  assign memOutput_0 = _zz_memInst_0_port0;
  assign _zz_memOutput_1 = io_fullRound;
  assign memOutput_1 = _zz_memInst_1_port0;
  assign _zz_memOutput_2 = io_fullRound;
  assign memOutput_2 = _zz_memInst_2_port0;
  assign _zz_memOutput_3 = io_fullRound;
  assign memOutput_3 = _zz_memInst_3_port0;
  assign _zz_memOutput_4 = io_fullRound;
  assign memOutput_4 = _zz_memInst_4_port0;
  assign _zz_memOutput_5 = io_fullRound;
  assign memOutput_5 = _zz_memInst_5_port0;
  assign _zz_memOutput_6 = io_fullRound;
  assign memOutput_6 = _zz_memInst_6_port0;
  assign _zz_memOutput_7 = io_fullRound;
  assign memOutput_7 = _zz_memInst_7_port0;
  assign _zz_memOutput_8 = io_fullRound;
  assign memOutput_8 = _zz_memInst_8_port0;
  assign _zz_memOutput_9 = io_fullRound;
  assign memOutput_9 = _zz_memInst_9_port0;
  assign _zz_memOutput_10 = io_fullRound;
  assign memOutput_10 = _zz_memInst_10_port0;
  assign _zz_memOutput_11 = io_fullRound;
  assign memOutput_11 = _zz_memInst_11_port0;
  assign io_constant = _zz_io_constant;

endmodule

module FullRoundConstantMem_2 (
  input      [3:0]    io_stateIndex,
  input      [2:0]    io_fullRound,
  output     [254:0]  io_constant
);

  wire       [254:0]  _zz_memInst_0_port0;
  wire       [254:0]  _zz_memInst_1_port0;
  wire       [254:0]  _zz_memInst_2_port0;
  wire       [254:0]  _zz_memInst_3_port0;
  wire       [254:0]  _zz_memInst_4_port0;
  wire       [254:0]  _zz_memInst_5_port0;
  wire       [254:0]  _zz_memInst_6_port0;
  wire       [254:0]  _zz_memInst_7_port0;
  wire       [254:0]  _zz_memInst_8_port0;
  reg        [254:0]  _zz_io_constant;
  wire       [253:0]  constantsMat_0_0;
  wire       [254:0]  constantsMat_0_1;
  wire       [254:0]  constantsMat_0_2;
  wire       [251:0]  constantsMat_0_3;
  wire       [251:0]  constantsMat_0_4;
  wire       [252:0]  constantsMat_0_5;
  wire       [253:0]  constantsMat_0_6;
  wire       [254:0]  constantsMat_0_7;
  wire       [254:0]  constantsMat_0_8;
  wire       [254:0]  constantsMat_1_0;
  wire       [247:0]  constantsMat_1_1;
  wire       [253:0]  constantsMat_1_2;
  wire       [252:0]  constantsMat_1_3;
  wire       [254:0]  constantsMat_1_4;
  wire       [254:0]  constantsMat_1_5;
  wire       [252:0]  constantsMat_1_6;
  wire       [253:0]  constantsMat_1_7;
  wire       [253:0]  constantsMat_1_8;
  wire       [253:0]  constantsMat_2_0;
  wire       [253:0]  constantsMat_2_1;
  wire       [254:0]  constantsMat_2_2;
  wire       [250:0]  constantsMat_2_3;
  wire       [251:0]  constantsMat_2_4;
  wire       [251:0]  constantsMat_2_5;
  wire       [253:0]  constantsMat_2_6;
  wire       [249:0]  constantsMat_2_7;
  wire       [254:0]  constantsMat_2_8;
  wire       [252:0]  constantsMat_3_0;
  wire       [253:0]  constantsMat_3_1;
  wire       [253:0]  constantsMat_3_2;
  wire       [254:0]  constantsMat_3_3;
  wire       [252:0]  constantsMat_3_4;
  wire       [253:0]  constantsMat_3_5;
  wire       [254:0]  constantsMat_3_6;
  wire       [254:0]  constantsMat_3_7;
  wire       [254:0]  constantsMat_3_8;
  wire       [254:0]  constantsMat_4_0;
  wire       [254:0]  constantsMat_4_1;
  wire       [253:0]  constantsMat_4_2;
  wire       [253:0]  constantsMat_4_3;
  wire       [254:0]  constantsMat_4_4;
  wire       [253:0]  constantsMat_4_5;
  wire       [250:0]  constantsMat_4_6;
  wire       [254:0]  constantsMat_4_7;
  wire       [254:0]  constantsMat_4_8;
  wire       [252:0]  constantsMat_5_0;
  wire       [251:0]  constantsMat_5_1;
  wire       [253:0]  constantsMat_5_2;
  wire       [254:0]  constantsMat_5_3;
  wire       [253:0]  constantsMat_5_4;
  wire       [253:0]  constantsMat_5_5;
  wire       [251:0]  constantsMat_5_6;
  wire       [254:0]  constantsMat_5_7;
  wire       [254:0]  constantsMat_5_8;
  wire       [252:0]  constantsMat_6_0;
  wire       [254:0]  constantsMat_6_1;
  wire       [253:0]  constantsMat_6_2;
  wire       [252:0]  constantsMat_6_3;
  wire       [251:0]  constantsMat_6_4;
  wire       [251:0]  constantsMat_6_5;
  wire       [253:0]  constantsMat_6_6;
  wire       [254:0]  constantsMat_6_7;
  wire       [254:0]  constantsMat_6_8;
  wire       [2:0]    _zz_memOutput_0;
  wire       [254:0]  memOutput_0;
  wire       [2:0]    _zz_memOutput_1;
  wire       [254:0]  memOutput_1;
  wire       [2:0]    _zz_memOutput_2;
  wire       [254:0]  memOutput_2;
  wire       [2:0]    _zz_memOutput_3;
  wire       [254:0]  memOutput_3;
  wire       [2:0]    _zz_memOutput_4;
  wire       [254:0]  memOutput_4;
  wire       [2:0]    _zz_memOutput_5;
  wire       [254:0]  memOutput_5;
  wire       [2:0]    _zz_memOutput_6;
  wire       [254:0]  memOutput_6;
  wire       [2:0]    _zz_memOutput_7;
  wire       [254:0]  memOutput_7;
  wire       [2:0]    _zz_memOutput_8;
  wire       [254:0]  memOutput_8;
  (* ram_style = "distributed" *) reg [254:0] memInst_0 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_1 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_2 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_3 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_4 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_5 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_6 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_7 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_8 [0:7];

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_6_memInst_0.bin",memInst_0);
  end
  assign _zz_memInst_0_port0 = memInst_0[_zz_memOutput_0];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_6_memInst_1.bin",memInst_1);
  end
  assign _zz_memInst_1_port0 = memInst_1[_zz_memOutput_1];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_6_memInst_2.bin",memInst_2);
  end
  assign _zz_memInst_2_port0 = memInst_2[_zz_memOutput_2];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_6_memInst_3.bin",memInst_3);
  end
  assign _zz_memInst_3_port0 = memInst_3[_zz_memOutput_3];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_6_memInst_4.bin",memInst_4);
  end
  assign _zz_memInst_4_port0 = memInst_4[_zz_memOutput_4];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_6_memInst_5.bin",memInst_5);
  end
  assign _zz_memInst_5_port0 = memInst_5[_zz_memOutput_5];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_6_memInst_6.bin",memInst_6);
  end
  assign _zz_memInst_6_port0 = memInst_6[_zz_memOutput_6];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_6_memInst_7.bin",memInst_7);
  end
  assign _zz_memInst_7_port0 = memInst_7[_zz_memOutput_7];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_6_memInst_8.bin",memInst_8);
  end
  assign _zz_memInst_8_port0 = memInst_8[_zz_memOutput_8];
  always @(*) begin
    case(io_stateIndex)
      4'b0000 : _zz_io_constant = memOutput_0;
      4'b0001 : _zz_io_constant = memOutput_1;
      4'b0010 : _zz_io_constant = memOutput_2;
      4'b0011 : _zz_io_constant = memOutput_3;
      4'b0100 : _zz_io_constant = memOutput_4;
      4'b0101 : _zz_io_constant = memOutput_5;
      4'b0110 : _zz_io_constant = memOutput_6;
      4'b0111 : _zz_io_constant = memOutput_7;
      default : _zz_io_constant = memOutput_8;
    endcase
  end

  assign constantsMat_0_0 = 254'h3e91e4318b42b3b46ab2eaa20758f1b7ce3e1b6e52db22a3bc9f62a154e12591;
  assign constantsMat_0_1 = 255'h606d462411d9478f9a64ef40a684bb8c9884df0a6d19f6c92148ea032ffdc233;
  assign constantsMat_0_2 = 255'h70eb12024b5286b643f1c0428aee5dcbefd428b6ade9f6fb95a876f3680e7895;
  assign constantsMat_0_3 = 252'hd30cc3ebc7c17a8c6536fa8ee214091f4a180242a4c6023991c8af69567a68d;
  assign constantsMat_0_4 = 252'h8de3def02284ee00844d5d83118fd29e7b6827a70b932217d0886604df13069;
  assign constantsMat_0_5 = 253'h18d50b44abaa91a94def29011b6cc16fd650c3a56841497949b0230afa0eb501;
  assign constantsMat_0_6 = 254'h2cab4d3bdb7e584a29d9ab5ab2b0677b3173fada1f689c626e7c9512adfebe3b;
  assign constantsMat_0_7 = 255'h696fb453b14ace8afeb635ebdbc8a5e4f003cdaf26729df803e875b077092734;
  assign constantsMat_0_8 = 255'h595b93471fd52b947757ad56e868f7d279dc3ba5137591a0dd1d87f1395d3e62;
  assign constantsMat_1_0 = 255'h5c066a52cbbf7e9e931eb4dee68cc07fe7ea951b3ef3f7f4e99f9eaf77b5a3fd;
  assign constantsMat_1_1 = 248'h8f48fc3455981bdc9b1a15445b53ee7803bd1db8ea54b91000e3c6d9749fa9;
  assign constantsMat_1_2 = 254'h27966b14eff60460a0c680b3e99fa04838dfd1c0df7974fc1f9dfa785b6d4c7b;
  assign constantsMat_1_3 = 253'h1af47a79ae038ba379c4930318059936721258e8768953c75f9be50188181ef3;
  assign constantsMat_1_4 = 255'h4da60fa08343a80d1d10358b1a842516c4a002e3213a1fd68da982fc706dfdd0;
  assign constantsMat_1_5 = 255'h506ce479f6829b116c531bb8701e60a30093f6e28152c665c2e7bb93e7f909c7;
  assign constantsMat_1_6 = 253'h1409146d455d78b5e6e772b8082b042c60e27cf27da8154ad2aad2b4bd9036d9;
  assign constantsMat_1_7 = 254'h3f358a561d88c192c47e12fae437fc71f1ed19f1ccfea988ea2cf6eaed45444e;
  assign constantsMat_1_8 = 254'h2c7e1bfc3a80b1d995169aaf03338c7f5df4a549c245105049b61964de5caa30;
  assign constantsMat_2_0 = 254'h3d22e0cb85842340ad544d9583f88c5a6802ef2901b79f329430e68add66283d;
  assign constantsMat_2_1 = 254'h367fb385b4abe7edb4d57662b4b61c55d0834825e1268b819e0b7d52808cdccc;
  assign constantsMat_2_2 = 255'h66b7ca7d5b7f35b888a7bf9d340a5bd7fba59f0ad626f76cb9578fcd99a56df3;
  assign constantsMat_2_3 = 251'h6f263dce27d7a44b526c21f14e49e3af42bd465562f92121f3ada8bfa36b105;
  assign constantsMat_2_4 = 252'h8b4e9fd2de81c5c21b5cfdc26c8efb4962f912ee7b31fe0ec242d3616058fa5;
  assign constantsMat_2_5 = 252'hd597246e65a88e1d7a3a08b611723476465c3826ca7272b96dadf217d7dfa91;
  assign constantsMat_2_6 = 254'h3c47484b1820082e4e033e3e2ff6fb4dab41da4a302303ba417960f2dbbd6309;
  assign constantsMat_2_7 = 250'h3bab48054d6906dbdbb52fbc44c61ae6bc487f3cf203e48d3c4022d47dca90e;
  assign constantsMat_2_8 = 255'h61aa65320ac4faa6002b4f5ab6b45c42606c06f345d6f9d354bb331e673addb6;
  assign constantsMat_3_0 = 253'h1985bf66cb7fc3b565a6f70c10c2e993209cf2a88cd5da50731597f22aeab17d;
  assign constantsMat_3_1 = 254'h30af9e128963614004f80e2900a40bc59c6ad722ea2ce15721b5c8914fdd1bd9;
  assign constantsMat_3_2 = 254'h2998a04579966d7ace93432b8fbe1d92f2821a10c69d382057346bd1c290c99f;
  assign constantsMat_3_3 = 255'h7185a2e4777cd0bbb325d04c94a9987ae9a43f1c901ac8d07e60d36ebf64b257;
  assign constantsMat_3_4 = 253'h1bd9efd9c6041cdbc3dbe928d1b8ed64dfdc54b8b60ef1aaf41338cf162f0b66;
  assign constantsMat_3_5 = 254'h25da6170bbf59cb09d42f191fddfa3f78cdeb7c822d7b0db2b3b698337c7db7a;
  assign constantsMat_3_6 = 255'h5ce067922bc0efb21f2e3bc6445da5d539a8912a6f0fbd2a92a4f4b219c90a95;
  assign constantsMat_3_7 = 255'h5f2a25117d18a8fd1e0ef4a3228cbbd554d71f907b26535efefff05b84bad092;
  assign constantsMat_3_8 = 255'h500e471d5259fa9f935120b4a4959aa9dad5c2b756a378a36ac4f4be35b5cb99;
  assign constantsMat_4_0 = 255'h63e5cf66ff63c50a7cc1142448d3c964919693ce9a0acff094163128944eff33;
  assign constantsMat_4_1 = 255'h53b1d3e06de9cd742c7a0e6c9006caadfd06ed13966af689a1d7c321b6a00404;
  assign constantsMat_4_2 = 254'h37bc7a0f8d588eb98fb98751355dc9376046b2c6833bf32755916eca9640fcf3;
  assign constantsMat_4_3 = 254'h3160b3e84a481a79866c183f6f58972a31d4b2656264fb5afbf6bdfb3323e7ac;
  assign constantsMat_4_4 = 255'h7377609f48b9505b08777ab52321b6dc6444aa93c911495f4dd1b10070a5cd9b;
  assign constantsMat_4_5 = 254'h2543fa7316becb685b6f1cb2233a666c26e7bba18d3f27e63a8b187865e4adbc;
  assign constantsMat_4_6 = 251'h6474819fd0ed10871680d953d068694b66548d8ec77993bb8abc56f7dc8cb90;
  assign constantsMat_4_7 = 255'h64db885dfdb21cf4d365f869d355ca1ed4b00d35bfb34807cf6421149a6130c0;
  assign constantsMat_4_8 = 255'h4f4784bf53e0185e61470da658ddc8a2a517bbd7771d8158d02aae8f5b740144;
  assign constantsMat_5_0 = 253'h1e09ce8cc4eded9d733d6cca1689b6dc18b659f22162fbd95232937754a517b1;
  assign constantsMat_5_1 = 252'habab92ef1505352dfe1475b832820eb0b4261c6b717dc942cef64771fb7b012;
  assign constantsMat_5_2 = 254'h2a456d5651e11c1e945eecb577f15b838077d892c177d9bc93057728d1476c4b;
  assign constantsMat_5_3 = 255'h5bc97ca566cb4bc80bc2621fe4c1f1b8ad4933736368ccfac5d5b3d90d40b1fc;
  assign constantsMat_5_4 = 254'h298eae333f5fcfb6951e8a1d84a538f683b29bd8366af001abd20cd0c1ab47dc;
  assign constantsMat_5_5 = 254'h2a37725bc58ffc48d9abefcd364737933659d44161112a920ca3459bea2a03af;
  assign constantsMat_5_6 = 252'he2180b1d5ab7d2742bc74f356713968de92ce656f427768b2c5f22275e9d877;
  assign constantsMat_5_7 = 255'h444aa434b1d479c486dda89b98162b7ccf461827ee8375d939fd575b95dbfaa9;
  assign constantsMat_5_8 = 255'h4421dc95a9cec1b543a5de52bbd000eaa78e1d5895ec875bcb00a746b8f3b544;
  assign constantsMat_6_0 = 253'h14ad89f435b3760ff99df873b6c649c9e861a288679a0b1fcbe329f4c6df8f03;
  assign constantsMat_6_1 = 255'h68e98d6b23b7f565c4e3944652eb0f6ec313bb5a6fa24a96cf8448c2ff3c981f;
  assign constantsMat_6_2 = 254'h34769b7079cc12b6e31b9090f2e1a250440493e4b10873142d0bfa591681b363;
  assign constantsMat_6_3 = 253'h1da019de812c83c3cc2f116bb9cd4f196618e69387bf881d573fe75dae84b4b6;
  assign constantsMat_6_4 = 252'ha4627715e3b5a550d2838528e443535ca8f7e75128fb470c60cace77afb03f2;
  assign constantsMat_6_5 = 252'hfb03b4a9106d2a8dc060de4fe4b6c8cc61dabcbce63b4d17ab92265b4371cb7;
  assign constantsMat_6_6 = 254'h239b18c7ad235b58a5324de832c492f43a327b0dc89d1c34ea715bd2aa94cf3e;
  assign constantsMat_6_7 = 255'h4bcdc12dc28664bad74f0cc5e28d8a1547a16a120d954241ee1cfc231e983474;
  assign constantsMat_6_8 = 255'h462a2815f18646d0d8958e2331ee6e19637b60314aba89a6b2a282e8d7ccef49;
  assign _zz_memOutput_0 = io_fullRound;
  assign memOutput_0 = _zz_memInst_0_port0;
  assign _zz_memOutput_1 = io_fullRound;
  assign memOutput_1 = _zz_memInst_1_port0;
  assign _zz_memOutput_2 = io_fullRound;
  assign memOutput_2 = _zz_memInst_2_port0;
  assign _zz_memOutput_3 = io_fullRound;
  assign memOutput_3 = _zz_memInst_3_port0;
  assign _zz_memOutput_4 = io_fullRound;
  assign memOutput_4 = _zz_memInst_4_port0;
  assign _zz_memOutput_5 = io_fullRound;
  assign memOutput_5 = _zz_memInst_5_port0;
  assign _zz_memOutput_6 = io_fullRound;
  assign memOutput_6 = _zz_memInst_6_port0;
  assign _zz_memOutput_7 = io_fullRound;
  assign memOutput_7 = _zz_memInst_7_port0;
  assign _zz_memOutput_8 = io_fullRound;
  assign memOutput_8 = _zz_memInst_8_port0;
  assign io_constant = _zz_io_constant;

endmodule

module FullRoundConstantMem_1 (
  input      [3:0]    io_stateIndex,
  input      [2:0]    io_fullRound,
  output     [254:0]  io_constant
);

  wire       [254:0]  _zz_memInst_0_port0;
  wire       [254:0]  _zz_memInst_1_port0;
  wire       [254:0]  _zz_memInst_2_port0;
  wire       [254:0]  _zz_memInst_3_port0;
  wire       [254:0]  _zz_memInst_4_port0;
  reg        [254:0]  _zz_io_constant;
  wire       [2:0]    _zz_io_constant_1;
  wire       [253:0]  constantsMat_0_0;
  wire       [254:0]  constantsMat_0_1;
  wire       [254:0]  constantsMat_0_2;
  wire       [254:0]  constantsMat_0_3;
  wire       [254:0]  constantsMat_0_4;
  wire       [254:0]  constantsMat_1_0;
  wire       [251:0]  constantsMat_1_1;
  wire       [249:0]  constantsMat_1_2;
  wire       [253:0]  constantsMat_1_3;
  wire       [254:0]  constantsMat_1_4;
  wire       [253:0]  constantsMat_2_0;
  wire       [253:0]  constantsMat_2_1;
  wire       [254:0]  constantsMat_2_2;
  wire       [253:0]  constantsMat_2_3;
  wire       [251:0]  constantsMat_2_4;
  wire       [253:0]  constantsMat_3_0;
  wire       [254:0]  constantsMat_3_1;
  wire       [254:0]  constantsMat_3_2;
  wire       [254:0]  constantsMat_3_3;
  wire       [253:0]  constantsMat_3_4;
  wire       [250:0]  constantsMat_4_0;
  wire       [251:0]  constantsMat_4_1;
  wire       [253:0]  constantsMat_4_2;
  wire       [254:0]  constantsMat_4_3;
  wire       [254:0]  constantsMat_4_4;
  wire       [254:0]  constantsMat_5_0;
  wire       [253:0]  constantsMat_5_1;
  wire       [254:0]  constantsMat_5_2;
  wire       [253:0]  constantsMat_5_3;
  wire       [254:0]  constantsMat_5_4;
  wire       [252:0]  constantsMat_6_0;
  wire       [254:0]  constantsMat_6_1;
  wire       [254:0]  constantsMat_6_2;
  wire       [254:0]  constantsMat_6_3;
  wire       [254:0]  constantsMat_6_4;
  wire       [2:0]    _zz_memOutput_0;
  wire       [254:0]  memOutput_0;
  wire       [2:0]    _zz_memOutput_1;
  wire       [254:0]  memOutput_1;
  wire       [2:0]    _zz_memOutput_2;
  wire       [254:0]  memOutput_2;
  wire       [2:0]    _zz_memOutput_3;
  wire       [254:0]  memOutput_3;
  wire       [2:0]    _zz_memOutput_4;
  wire       [254:0]  memOutput_4;
  (* ram_style = "distributed" *) reg [254:0] memInst_0 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_1 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_2 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_3 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_4 [0:7];

  assign _zz_io_constant_1 = io_stateIndex[2:0];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_5_memInst_0.bin",memInst_0);
  end
  assign _zz_memInst_0_port0 = memInst_0[_zz_memOutput_0];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_5_memInst_1.bin",memInst_1);
  end
  assign _zz_memInst_1_port0 = memInst_1[_zz_memOutput_1];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_5_memInst_2.bin",memInst_2);
  end
  assign _zz_memInst_2_port0 = memInst_2[_zz_memOutput_2];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_5_memInst_3.bin",memInst_3);
  end
  assign _zz_memInst_3_port0 = memInst_3[_zz_memOutput_3];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_5_memInst_4.bin",memInst_4);
  end
  assign _zz_memInst_4_port0 = memInst_4[_zz_memOutput_4];
  always @(*) begin
    case(_zz_io_constant_1)
      3'b000 : _zz_io_constant = memOutput_0;
      3'b001 : _zz_io_constant = memOutput_1;
      3'b010 : _zz_io_constant = memOutput_2;
      3'b011 : _zz_io_constant = memOutput_3;
      default : _zz_io_constant = memOutput_4;
    endcase
  end

  assign constantsMat_0_0 = 254'h3e90d6cd6c7833beea8072690272c364efb62462b729ba3562df178936cee858;
  assign constantsMat_0_1 = 255'h5b15a4cbaf84cb6230e39b5b4a7430dc05d6d9b02812267bb2bfa42f73df7ae2;
  assign constantsMat_0_2 = 255'h58ca12da49ef4ab21f950964eae842a1970bf09ebf6d1b94d4933b1b4e728ee9;
  assign constantsMat_0_3 = 255'h7290a0e823d4fdc123c122b2e0abddf01ec1af883fe512210beaa100831b5c1c;
  assign constantsMat_0_4 = 255'h49356536fd1d9842465dabd0935b9703d5c3d9009dc1c9b30cc2836ed64f4ad0;
  assign constantsMat_1_0 = 255'h6253f8445181947e7ce6886a71222e22c791d2fe42433fad63f21b32a6d4c501;
  assign constantsMat_1_1 = 252'hb0a1c20e1a89b10db06e7c3d5536dfe9cf13e57c92ee940943c1f285ac1c66f;
  assign constantsMat_1_2 = 250'h2d70f909d350eb69e1ae4db73c91d81bf2327b62f54b6a11a57147d9c209055;
  assign constantsMat_1_3 = 254'h2a8b5c7582103c71bc617b5161fc3ff2d686f36f8b4115c9725bbf69e3f6bd6a;
  assign constantsMat_1_4 = 255'h717b04c11072646d75a9ea620113af3a34b44f37ded6f065effeb9206e4114ed;
  assign constantsMat_2_0 = 254'h39102cfe4976829c17350bef3ce413f7090a1d1f8dd915bf0029823895b6df77;
  assign constantsMat_2_1 = 254'h268f30e1d558361ef8e6a425541a6d224870ba6e333f13efbe3d9f908da0aa79;
  assign constantsMat_2_2 = 255'h41878a1395ae763c0db29b1a3fd1a0b8632a6665db7298bc7d09b9ec9134abe2;
  assign constantsMat_2_3 = 254'h30c09edc44a3b6fc25dc04c842aea1849f39a71449a1549c3508eed65cb2af91;
  assign constantsMat_2_4 = 252'hdd2e613dfddf86a22c821832a867d87eedd40f4aca1a1ff463c03b14fda248e;
  assign constantsMat_3_0 = 254'h34f0bc9689c7a8bfdcfd4a28bb3591b062b9fb610571b4e77183603603c824f3;
  assign constantsMat_3_1 = 255'h637ba50bbf8f4cbc618ae65d2ee1314dce4528feb68cf0e96f258cec4753f58f;
  assign constantsMat_3_2 = 255'h52188f75db41ed39d3d8775d2cf76ecea4657029d1b18211075c49ae16f0b559;
  assign constantsMat_3_3 = 255'h6eef08529ac5126c3c0456985fadaee5dd169a00fd55409a0051f1fad894717e;
  assign constantsMat_3_4 = 254'h2be380692474498fb20d6c8ed7eb94a693faf8b6f80cbd0cb82526c6857c31af;
  assign constantsMat_4_0 = 251'h56d28c7bdc6b5c23534e8c14987ebeb834add7427ded651c69dc23e27120456;
  assign constantsMat_4_1 = 252'hcb487276eced6a6e144ac2b4a17a00bbae913c586008f1a3c762c83fc588e6e;
  assign constantsMat_4_2 = 254'h35a019c05a9ed06b228da72f5305348809401a868b0089f32c7718717c7a50a8;
  assign constantsMat_4_3 = 255'h711af051b3f23397c815a0554d315eae13fbddbfb38a14704201eccfb2506a6a;
  assign constantsMat_4_4 = 255'h692fbd6f78cc46ad074223fe12c2e188d6270453a760e7b2210701ae5cb0a954;
  assign constantsMat_5_0 = 255'h54fff081f436a8125535858ccbee9f056fcfc9c27345b28680ee08141584ac15;
  assign constantsMat_5_1 = 254'h307faf11551f916c049b8b283d6d0f5dd0576d3c2d22b95c7e68dbc5056c2ca0;
  assign constantsMat_5_2 = 255'h618a5d16dd4c250c185682b1dc0177c19a8dc18fd5d55bf001c674dfefa067a4;
  assign constantsMat_5_3 = 254'h240cbef05002149467cd0286e8b919db13f7abeb261359957170dc3e83a591b0;
  assign constantsMat_5_4 = 255'h5b5e10efc9f91a8b417bc7de959d984f5906efe76291c3d11c52c684668fce23;
  assign constantsMat_6_0 = 253'h1e02df65cba9f57559f54e595e8e1b929538b86c1f93f66fabb318eb21854b3b;
  assign constantsMat_6_1 = 255'h4ef39debb5bcc97c9a3e4453ec20d7e83df165527d82d032fc161bb46f046958;
  assign constantsMat_6_2 = 255'h6ca2cb9e63ceab96e58eb55a293080b16e037935448d7f83d65ce0841fb1f453;
  assign constantsMat_6_3 = 255'h5d466700cccb3c5415d47a795b146ce17634043fffecedc55952e9ec80c4d3ac;
  assign constantsMat_6_4 = 255'h65e2e8377190483bc6c095638c9fcce83369f3454fba50fbc37cab22808060ce;
  assign _zz_memOutput_0 = io_fullRound;
  assign memOutput_0 = _zz_memInst_0_port0;
  assign _zz_memOutput_1 = io_fullRound;
  assign memOutput_1 = _zz_memInst_1_port0;
  assign _zz_memOutput_2 = io_fullRound;
  assign memOutput_2 = _zz_memInst_2_port0;
  assign _zz_memOutput_3 = io_fullRound;
  assign memOutput_3 = _zz_memInst_3_port0;
  assign _zz_memOutput_4 = io_fullRound;
  assign memOutput_4 = _zz_memInst_4_port0;
  assign io_constant = _zz_io_constant;

endmodule

module FullRoundConstantMem (
  input      [3:0]    io_stateIndex,
  input      [2:0]    io_fullRound,
  output     [254:0]  io_constant
);

  wire       [254:0]  _zz_memInst_0_port0;
  wire       [254:0]  _zz_memInst_1_port0;
  wire       [254:0]  _zz_memInst_2_port0;
  reg        [254:0]  _zz_io_constant;
  wire       [1:0]    _zz_io_constant_1;
  wire       [254:0]  constantsMat_0_0;
  wire       [253:0]  constantsMat_0_1;
  wire       [253:0]  constantsMat_0_2;
  wire       [254:0]  constantsMat_1_0;
  wire       [254:0]  constantsMat_1_1;
  wire       [254:0]  constantsMat_1_2;
  wire       [249:0]  constantsMat_2_0;
  wire       [254:0]  constantsMat_2_1;
  wire       [254:0]  constantsMat_2_2;
  wire       [252:0]  constantsMat_3_0;
  wire       [253:0]  constantsMat_3_1;
  wire       [254:0]  constantsMat_3_2;
  wire       [254:0]  constantsMat_4_0;
  wire       [252:0]  constantsMat_4_1;
  wire       [253:0]  constantsMat_4_2;
  wire       [254:0]  constantsMat_5_0;
  wire       [253:0]  constantsMat_5_1;
  wire       [253:0]  constantsMat_5_2;
  wire       [253:0]  constantsMat_6_0;
  wire       [254:0]  constantsMat_6_1;
  wire       [254:0]  constantsMat_6_2;
  wire       [2:0]    _zz_memOutput_0;
  wire       [254:0]  memOutput_0;
  wire       [2:0]    _zz_memOutput_1;
  wire       [254:0]  memOutput_1;
  wire       [2:0]    _zz_memOutput_2;
  wire       [254:0]  memOutput_2;
  (* ram_style = "distributed" *) reg [254:0] memInst_0 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_1 [0:7];
  (* ram_style = "distributed" *) reg [254:0] memInst_2 [0:7];

  assign _zz_io_constant_1 = io_stateIndex[1:0];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_4_memInst_0.bin",memInst_0);
  end
  assign _zz_memInst_0_port0 = memInst_0[_zz_memOutput_0];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_4_memInst_1.bin",memInst_1);
  end
  assign _zz_memInst_1_port0 = memInst_1[_zz_memOutput_1];
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_AddRoundConstantStage_constantMemory_fullRoundConstantMem_4_memInst_2.bin",memInst_2);
  end
  assign _zz_memInst_2_port0 = memInst_2[_zz_memOutput_2];
  always @(*) begin
    case(_zz_io_constant_1)
      2'b00 : _zz_io_constant = memOutput_0;
      2'b01 : _zz_io_constant = memOutput_1;
      default : _zz_io_constant = memOutput_2;
    endcase
  end

  assign constantsMat_0_0 = 255'h4517ba4b7c09e98c9f5655bc5716a24850897887d3a35419f94ac1947de7dfbf;
  assign constantsMat_0_1 = 254'h2924588522082c34139f0c1aa9387186f70629ecb6bc61c8634c4c5d1e922f65;
  assign constantsMat_0_2 = 254'h2176e2a8e17b0334d1a9afd2c536e7c1f53c66223285900202e3da796b2588e7;
  assign constantsMat_1_0 = 255'h59007dc06b70d92913d9f5410992584bd22848ff29a3a26a3357a3e5fb0e2c83;
  assign constantsMat_1_1 = 255'h49855421a67d44da22ca7e6753629da1de5f847ccbb3bcecba279ba13e25d236;
  assign constantsMat_1_2 = 255'h4cc12f94e93b10143c09313a651e91f1e8e91b06e0f3c15a36bc60adb18fb495;
  assign constantsMat_2_0 = 250'h36cd8b4d3835fc3d14da6d2cb573ee6b78f297c66af464f8ae4508d9adf8c1c;
  assign constantsMat_2_1 = 255'h72a2a116737f0d1b362f024b68a823d31070dabe5f80fcd95b7c05b57a4a9bbd;
  assign constantsMat_2_2 = 255'h577c0b4f62187b7d212d7faafaba0cd3bde34183bbdcc676307734828b5f8720;
  assign constantsMat_3_0 = 253'h1cb041121f1c945cc101ff983bc06262946b768466e29527b7c615ac86a51179;
  assign constantsMat_3_1 = 254'h2799270041b61254b3e55fc6376c34c22babe8e7aefca45941bbd60571403aa8;
  assign constantsMat_3_2 = 255'h548c7c2ab82f5dc355c98968cb3faddc2ce697691ec4afd772191dd45f75f510;
  assign constantsMat_4_0 = 255'h56c50a0987544b0ae2cebf0f4ffc771e378a357925dbe02f121a624ff2fa6515;
  assign constantsMat_4_1 = 253'h1c9b4c2f0347c4380a9ce5dbdff12dea75796d32e375f949eef3d92cdb1a75de;
  assign constantsMat_4_2 = 254'h3ae634d0aee1b659a7a5fe04ba22cfe642118279e686b956a43fce9c67ff43e2;
  assign constantsMat_5_0 = 255'h4e3f7b301f96c62eae42227521870e8676c24cf7ff4dc0a2f6250e0e77939021;
  assign constantsMat_5_1 = 254'h32027f4b29ba5dfa718a63356b649250792599b022051241e04b4510e65a7396;
  assign constantsMat_5_2 = 254'h24487f8a7ac6a8c44795688b5d429175192d25e5d172fcda75865a2e698aa5e0;
  assign constantsMat_6_0 = 254'h2698a559226880614d3fe274a97b265f43f6e6aae098b314b6548061f3d6d4a2;
  assign constantsMat_6_1 = 255'h697c358044a0ea98cdc5e04faf0acbc8deb7495a7c56cc6ffeb966f1ad59f50e;
  assign constantsMat_6_2 = 255'h5a9296c00ddd3f06b34412fe6a6cbea2fcb8abcd549d64cbae9ae8329d3ba5e5;
  assign _zz_memOutput_0 = io_fullRound;
  assign memOutput_0 = _zz_memInst_0_port0;
  assign _zz_memOutput_1 = io_fullRound;
  assign memOutput_1 = _zz_memInst_1_port0;
  assign _zz_memOutput_2 = io_fullRound;
  assign memOutput_2 = _zz_memInst_2_port0;
  assign io_constant = _zz_io_constant;

endmodule

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

//ShiftRegister replaced by ShiftRegister

module ShiftRegister (
  input               io_ena,
  input               io_init,
  input      [254:0]  io_serialInput,
  input      [254:0]  io_parallelInput_0,
  input      [254:0]  io_parallelInput_1,
  input      [254:0]  io_parallelInput_2,
  input      [254:0]  io_parallelInput_3,
  input      [254:0]  io_parallelInput_4,
  input      [254:0]  io_parallelInput_5,
  input      [254:0]  io_parallelInput_6,
  input      [254:0]  io_parallelInput_7,
  input      [254:0]  io_parallelInput_8,
  input      [254:0]  io_parallelInput_9,
  input      [254:0]  io_parallelInput_10,
  input      [254:0]  io_parallelInput_11,
  output     [254:0]  io_parallelOutput_0,
  output     [254:0]  io_parallelOutput_1,
  output     [254:0]  io_parallelOutput_2,
  output     [254:0]  io_parallelOutput_3,
  output     [254:0]  io_parallelOutput_4,
  output     [254:0]  io_parallelOutput_5,
  output     [254:0]  io_parallelOutput_6,
  output     [254:0]  io_parallelOutput_7,
  output     [254:0]  io_parallelOutput_8,
  output     [254:0]  io_parallelOutput_9,
  output     [254:0]  io_parallelOutput_10,
  output     [254:0]  io_parallelOutput_11,
  input               clk,
  input               resetn
);

  wire       [254:0]  _zz__zz_io_parallelOutput_0;
  wire       [254:0]  _zz__zz_io_parallelOutput_0_1;
  wire       [254:0]  _zz__zz_buffer_0;
  wire       [254:0]  _zz__zz_buffer_0_1;
  reg        [254:0]  buffer_0;
  reg        [254:0]  buffer_1;
  reg        [254:0]  buffer_2;
  reg        [254:0]  buffer_3;
  reg        [254:0]  buffer_4;
  reg        [254:0]  buffer_5;
  reg        [254:0]  buffer_6;
  reg        [254:0]  buffer_7;
  reg        [254:0]  buffer_8;
  reg        [254:0]  buffer_9;
  reg        [254:0]  buffer_10;
  reg        [254:0]  buffer_11;
  wire       [3059:0] _zz_io_parallelOutput_0;
  wire       [3059:0] _zz_buffer_0;

  assign _zz__zz_io_parallelOutput_0 = buffer_1;
  assign _zz__zz_io_parallelOutput_0_1 = buffer_0;
  assign _zz__zz_buffer_0 = io_parallelInput_1;
  assign _zz__zz_buffer_0_1 = io_parallelInput_0;
  assign _zz_io_parallelOutput_0 = {buffer_11,{buffer_10,{buffer_9,{buffer_8,{buffer_7,{buffer_6,{buffer_5,{buffer_4,{buffer_3,{buffer_2,{_zz__zz_io_parallelOutput_0,_zz__zz_io_parallelOutput_0_1}}}}}}}}}}};
  assign io_parallelOutput_0 = _zz_io_parallelOutput_0[254 : 0];
  assign io_parallelOutput_1 = _zz_io_parallelOutput_0[509 : 255];
  assign io_parallelOutput_2 = _zz_io_parallelOutput_0[764 : 510];
  assign io_parallelOutput_3 = _zz_io_parallelOutput_0[1019 : 765];
  assign io_parallelOutput_4 = _zz_io_parallelOutput_0[1274 : 1020];
  assign io_parallelOutput_5 = _zz_io_parallelOutput_0[1529 : 1275];
  assign io_parallelOutput_6 = _zz_io_parallelOutput_0[1784 : 1530];
  assign io_parallelOutput_7 = _zz_io_parallelOutput_0[2039 : 1785];
  assign io_parallelOutput_8 = _zz_io_parallelOutput_0[2294 : 2040];
  assign io_parallelOutput_9 = _zz_io_parallelOutput_0[2549 : 2295];
  assign io_parallelOutput_10 = _zz_io_parallelOutput_0[2804 : 2550];
  assign io_parallelOutput_11 = _zz_io_parallelOutput_0[3059 : 2805];
  assign _zz_buffer_0 = {io_parallelInput_11,{io_parallelInput_10,{io_parallelInput_9,{io_parallelInput_8,{io_parallelInput_7,{io_parallelInput_6,{io_parallelInput_5,{io_parallelInput_4,{io_parallelInput_3,{io_parallelInput_2,{_zz__zz_buffer_0,_zz__zz_buffer_0_1}}}}}}}}}}};
  always @(posedge clk) begin
    if(!resetn) begin
      buffer_0 <= 255'h0;
      buffer_1 <= 255'h0;
      buffer_2 <= 255'h0;
      buffer_3 <= 255'h0;
      buffer_4 <= 255'h0;
      buffer_5 <= 255'h0;
      buffer_6 <= 255'h0;
      buffer_7 <= 255'h0;
      buffer_8 <= 255'h0;
      buffer_9 <= 255'h0;
      buffer_10 <= 255'h0;
      buffer_11 <= 255'h0;
    end else begin
      if(io_init) begin
        buffer_0 <= _zz_buffer_0[254 : 0];
        buffer_1 <= _zz_buffer_0[509 : 255];
        buffer_2 <= _zz_buffer_0[764 : 510];
        buffer_3 <= _zz_buffer_0[1019 : 765];
        buffer_4 <= _zz_buffer_0[1274 : 1020];
        buffer_5 <= _zz_buffer_0[1529 : 1275];
        buffer_6 <= _zz_buffer_0[1784 : 1530];
        buffer_7 <= _zz_buffer_0[2039 : 1785];
        buffer_8 <= _zz_buffer_0[2294 : 2040];
        buffer_9 <= _zz_buffer_0[2549 : 2295];
        buffer_10 <= _zz_buffer_0[2804 : 2550];
        buffer_11 <= _zz_buffer_0[3059 : 2805];
      end else begin
        if(io_ena) begin
          buffer_0 <= io_serialInput;
          buffer_1 <= buffer_0;
          buffer_2 <= buffer_1;
          buffer_3 <= buffer_2;
          buffer_4 <= buffer_3;
          buffer_5 <= buffer_4;
          buffer_6 <= buffer_5;
          buffer_7 <= buffer_6;
          buffer_8 <= buffer_7;
          buffer_9 <= buffer_8;
          buffer_10 <= buffer_9;
          buffer_11 <= buffer_10;
        end
      end
    end
  end


endmodule

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

//ModAdderPiped replaced by ModAdderPiped

module ModAdderPiped (
  input      [254:0]  io_op1,
  input      [254:0]  io_op2,
  output     [254:0]  io_res,
  input               clk,
  input               resetn
);

  wire       [254:0]  simAdderIP_49_io_inputA;
  wire       [255:0]  simAdderIP_48_io_outputS;
  wire       [255:0]  simAdderIP_49_io_outputS;
  wire       [255:0]  _zz_io_res;
  reg        [255:0]  simAdderIP_48_io_outputS_delay_1;
  reg        [255:0]  simAdderIP_48_io_outputS_delay_2;
  reg        [255:0]  simAdderIP_48_io_outputS_delay_3;
  reg        [255:0]  simAdderIP_48_io_outputS_delay_4;
  reg        [255:0]  simAdderIP_48_io_outputS_delay_5;
  reg        [255:0]  simAdderIP_48_io_outputS_delay_6;
  reg        [255:0]  simAdderIP_48_io_outputS_delay_7;
  reg        [255:0]  adderRes1Delayed;

  assign _zz_io_res = ((adderRes1Delayed[255] || simAdderIP_49_io_outputS[255]) ? simAdderIP_49_io_outputS : adderRes1Delayed);
  SimAdderIP simAdderIP_48 (
    .io_inputA     (io_op1[254:0]                    ), //i
    .io_inputB     (io_op2[254:0]                    ), //i
    .io_outputS    (simAdderIP_48_io_outputS[255:0]  ), //o
    .clk           (clk                              ), //i
    .resetn        (resetn                           )  //i
  );
  SimAdderIP simAdderIP_49 (
    .io_inputA     (simAdderIP_49_io_inputA[254:0]                                         ), //i
    .io_inputB     (255'h0c1258acd66282b7ccc627f7f65e27faac425bfd0001a40100000000ffffffff  ), //i
    .io_outputS    (simAdderIP_49_io_outputS[255:0]                                        ), //o
    .clk           (clk                                                                    ), //i
    .resetn        (resetn                                                                 )  //i
  );
  assign simAdderIP_49_io_inputA = simAdderIP_48_io_outputS[254:0];
  assign io_res = _zz_io_res[254:0];
  always @(posedge clk) begin
    simAdderIP_48_io_outputS_delay_1 <= simAdderIP_48_io_outputS;
    simAdderIP_48_io_outputS_delay_2 <= simAdderIP_48_io_outputS_delay_1;
    simAdderIP_48_io_outputS_delay_3 <= simAdderIP_48_io_outputS_delay_2;
    simAdderIP_48_io_outputS_delay_4 <= simAdderIP_48_io_outputS_delay_3;
    simAdderIP_48_io_outputS_delay_5 <= simAdderIP_48_io_outputS_delay_4;
    simAdderIP_48_io_outputS_delay_6 <= simAdderIP_48_io_outputS_delay_5;
    simAdderIP_48_io_outputS_delay_7 <= simAdderIP_48_io_outputS_delay_6;
    adderRes1Delayed <= simAdderIP_48_io_outputS_delay_7;
  end


endmodule

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow_1 replaced by MultiplierFlow_1

//MultiplierFlow replaced by MultiplierFlow

//MultiplierFlow_1 replaced by MultiplierFlow_1

module MultiplierFlow_1 (
  input               io_input_valid,
  input      [255:0]  io_input_payload_op1,
  input      [255:0]  io_input_payload_op2,
  output              io_output_valid,
  output     [511:0]  io_output_payload_res,
  input               clk,
  input               resetn
);

  wire       [33:0]   multiplierIPFlow_1215_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1215_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1216_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1216_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1218_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1218_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1219_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1219_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1221_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1221_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1222_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1222_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1224_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1224_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1225_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1225_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1227_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1227_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1228_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1228_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1230_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1230_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1231_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1231_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1233_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1233_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1234_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1234_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1236_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1236_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1237_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1237_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1239_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1239_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1240_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1240_io_input_payload_op2;
  wire                multiplierIPFlow_1215_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1215_io_output_payload_res;
  wire                multiplierIPFlow_1216_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1216_io_output_payload_res;
  wire                multiplierIPFlow_1217_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1217_io_output_payload_res;
  wire                multiplierIPFlow_1218_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1218_io_output_payload_res;
  wire                multiplierIPFlow_1219_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1219_io_output_payload_res;
  wire                multiplierIPFlow_1220_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1220_io_output_payload_res;
  wire                multiplierIPFlow_1221_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1221_io_output_payload_res;
  wire                multiplierIPFlow_1222_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1222_io_output_payload_res;
  wire                multiplierIPFlow_1223_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1223_io_output_payload_res;
  wire                multiplierIPFlow_1224_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1224_io_output_payload_res;
  wire                multiplierIPFlow_1225_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1225_io_output_payload_res;
  wire                multiplierIPFlow_1226_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1226_io_output_payload_res;
  wire                multiplierIPFlow_1227_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1227_io_output_payload_res;
  wire                multiplierIPFlow_1228_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1228_io_output_payload_res;
  wire                multiplierIPFlow_1229_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1229_io_output_payload_res;
  wire                multiplierIPFlow_1230_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1230_io_output_payload_res;
  wire                multiplierIPFlow_1231_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1231_io_output_payload_res;
  wire                multiplierIPFlow_1232_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1232_io_output_payload_res;
  wire                multiplierIPFlow_1233_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1233_io_output_payload_res;
  wire                multiplierIPFlow_1234_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1234_io_output_payload_res;
  wire                multiplierIPFlow_1235_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1235_io_output_payload_res;
  wire                multiplierIPFlow_1236_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1236_io_output_payload_res;
  wire                multiplierIPFlow_1237_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1237_io_output_payload_res;
  wire                multiplierIPFlow_1238_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1238_io_output_payload_res;
  wire                multiplierIPFlow_1239_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1239_io_output_payload_res;
  wire                multiplierIPFlow_1240_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1240_io_output_payload_res;
  wire                multiplierIPFlow_1241_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1241_io_output_payload_res;
  wire       [65:0]   _zz__zz_io_input_payload_op1_10;
  wire       [64:0]   _zz__zz_io_input_payload_op1_10_1;
  wire       [65:0]   _zz__zz_io_input_payload_op2_10;
  wire       [64:0]   _zz__zz_io_input_payload_op2_10_1;
  wire       [67:0]   _zz__zz_output_payload_res_2;
  wire       [67:0]   _zz__zz_output_payload_res_2_1;
  wire       [131:0]  _zz__zz_output_payload_res_3;
  wire       [131:0]  _zz__zz_output_payload_res_3_1;
  wire       [131:0]  _zz__zz_output_payload_res_3_2;
  wire       [131:0]  _zz__zz_output_payload_res_3_3;
  wire       [99:0]   _zz__zz_output_payload_res_3_4;
  wire       [67:0]   _zz__zz_output_payload_res_6;
  wire       [67:0]   _zz__zz_output_payload_res_6_1;
  wire       [131:0]  _zz__zz_output_payload_res_7;
  wire       [131:0]  _zz__zz_output_payload_res_7_1;
  wire       [131:0]  _zz__zz_output_payload_res_7_2;
  wire       [131:0]  _zz__zz_output_payload_res_7_3;
  wire       [99:0]   _zz__zz_output_payload_res_7_4;
  wire       [67:0]   _zz__zz_output_payload_res_10;
  wire       [67:0]   _zz__zz_output_payload_res_10_1;
  wire       [131:0]  _zz__zz_output_payload_res_11;
  wire       [131:0]  _zz__zz_output_payload_res_11_1;
  wire       [131:0]  _zz__zz_output_payload_res_11_2;
  wire       [131:0]  _zz__zz_output_payload_res_11_3;
  wire       [99:0]   _zz__zz_output_payload_res_11_4;
  wire       [131:0]  _zz__zz_output_payload_res_14;
  wire       [131:0]  _zz__zz_output_payload_res_14_1;
  wire       [259:0]  _zz__zz_output_payload_res_15;
  wire       [259:0]  _zz__zz_output_payload_res_15_1;
  wire       [259:0]  _zz__zz_output_payload_res_15_2;
  wire       [259:0]  _zz__zz_output_payload_res_15_3;
  wire       [259:0]  _zz__zz_output_payload_res_15_4;
  wire       [195:0]  _zz__zz_output_payload_res_15_5;
  wire       [65:0]   _zz__zz_io_input_payload_op1_34;
  wire       [64:0]   _zz__zz_io_input_payload_op1_34_1;
  wire       [65:0]   _zz__zz_io_input_payload_op2_34;
  wire       [64:0]   _zz__zz_io_input_payload_op2_34_1;
  wire       [67:0]   _zz__zz_output_payload_res_18;
  wire       [67:0]   _zz__zz_output_payload_res_18_1;
  wire       [131:0]  _zz__zz_output_payload_res_19;
  wire       [131:0]  _zz__zz_output_payload_res_19_1;
  wire       [131:0]  _zz__zz_output_payload_res_19_2;
  wire       [131:0]  _zz__zz_output_payload_res_19_3;
  wire       [99:0]   _zz__zz_output_payload_res_19_4;
  wire       [67:0]   _zz__zz_output_payload_res_22;
  wire       [67:0]   _zz__zz_output_payload_res_22_1;
  wire       [131:0]  _zz__zz_output_payload_res_23;
  wire       [131:0]  _zz__zz_output_payload_res_23_1;
  wire       [131:0]  _zz__zz_output_payload_res_23_2;
  wire       [131:0]  _zz__zz_output_payload_res_23_3;
  wire       [99:0]   _zz__zz_output_payload_res_23_4;
  wire       [67:0]   _zz__zz_output_payload_res_26;
  wire       [67:0]   _zz__zz_output_payload_res_26_1;
  wire       [131:0]  _zz__zz_output_payload_res_27;
  wire       [131:0]  _zz__zz_output_payload_res_27_1;
  wire       [131:0]  _zz__zz_output_payload_res_27_2;
  wire       [131:0]  _zz__zz_output_payload_res_27_3;
  wire       [99:0]   _zz__zz_output_payload_res_27_4;
  wire       [131:0]  _zz__zz_output_payload_res_30;
  wire       [131:0]  _zz__zz_output_payload_res_30_1;
  wire       [259:0]  _zz__zz_output_payload_res_31;
  wire       [259:0]  _zz__zz_output_payload_res_31_1;
  wire       [259:0]  _zz__zz_output_payload_res_31_2;
  wire       [259:0]  _zz__zz_output_payload_res_31_3;
  wire       [259:0]  _zz__zz_output_payload_res_31_4;
  wire       [195:0]  _zz__zz_output_payload_res_31_5;
  wire       [65:0]   _zz__zz_io_input_payload_op1_58;
  wire       [64:0]   _zz__zz_io_input_payload_op1_58_1;
  wire       [65:0]   _zz__zz_io_input_payload_op2_58;
  wire       [64:0]   _zz__zz_io_input_payload_op2_58_1;
  wire       [67:0]   _zz__zz_output_payload_res_34;
  wire       [67:0]   _zz__zz_output_payload_res_34_1;
  wire       [131:0]  _zz__zz_output_payload_res_35;
  wire       [131:0]  _zz__zz_output_payload_res_35_1;
  wire       [131:0]  _zz__zz_output_payload_res_35_2;
  wire       [131:0]  _zz__zz_output_payload_res_35_3;
  wire       [99:0]   _zz__zz_output_payload_res_35_4;
  wire       [67:0]   _zz__zz_output_payload_res_38;
  wire       [67:0]   _zz__zz_output_payload_res_38_1;
  wire       [131:0]  _zz__zz_output_payload_res_39;
  wire       [131:0]  _zz__zz_output_payload_res_39_1;
  wire       [131:0]  _zz__zz_output_payload_res_39_2;
  wire       [131:0]  _zz__zz_output_payload_res_39_3;
  wire       [99:0]   _zz__zz_output_payload_res_39_4;
  wire       [67:0]   _zz__zz_output_payload_res_42;
  wire       [67:0]   _zz__zz_output_payload_res_42_1;
  wire       [131:0]  _zz__zz_output_payload_res_43;
  wire       [131:0]  _zz__zz_output_payload_res_43_1;
  wire       [131:0]  _zz__zz_output_payload_res_43_2;
  wire       [131:0]  _zz__zz_output_payload_res_43_3;
  wire       [99:0]   _zz__zz_output_payload_res_43_4;
  wire       [131:0]  _zz__zz_output_payload_res_46;
  wire       [131:0]  _zz__zz_output_payload_res_46_1;
  wire       [259:0]  _zz__zz_output_payload_res_47;
  wire       [259:0]  _zz__zz_output_payload_res_47_1;
  wire       [259:0]  _zz__zz_output_payload_res_47_2;
  wire       [259:0]  _zz__zz_output_payload_res_47_3;
  wire       [259:0]  _zz__zz_output_payload_res_47_4;
  wire       [195:0]  _zz__zz_output_payload_res_47_5;
  wire       [257:0]  _zz__zz_output_payload_res_50;
  wire       [257:0]  _zz__zz_output_payload_res_50_1;
  wire       [511:0]  _zz_output_payload_res_51;
  wire       [511:0]  _zz_output_payload_res_52;
  wire       [511:0]  _zz_output_payload_res_53;
  wire       [511:0]  _zz_output_payload_res_54;
  wire       [384:0]  _zz_output_payload_res_55;
  wire       [127:0]  _zz_io_input_payload_op1;
  wire       [127:0]  _zz_io_input_payload_op1_1;
  wire       [127:0]  _zz_io_input_payload_op2;
  wire       [127:0]  _zz_io_input_payload_op2_1;
  reg                 _zz_io_input_valid;
  reg        [127:0]  _zz_io_input_payload_op1_2;
  reg        [127:0]  _zz_io_input_payload_op1_3;
  reg        [127:0]  _zz_io_input_payload_op2_2;
  reg        [127:0]  _zz_io_input_payload_op2_3;
  reg        [128:0]  _zz_io_input_payload_op1_4;
  reg        [128:0]  _zz_io_input_payload_op2_4;
  wire       [128:0]  _zz_io_input_payload_op1_5;
  wire       [128:0]  _zz_io_input_payload_op2_5;
  wire       [64:0]   _zz_io_input_payload_op1_6;
  wire       [63:0]   _zz_io_input_payload_op1_7;
  wire       [64:0]   _zz_io_input_payload_op2_6;
  wire       [63:0]   _zz_io_input_payload_op2_7;
  reg                 _zz_io_input_valid_1;
  reg        [64:0]   _zz_io_input_payload_op1_8;
  reg        [63:0]   _zz_io_input_payload_op1_9;
  reg        [64:0]   _zz_io_input_payload_op2_8;
  reg        [63:0]   _zz_io_input_payload_op2_9;
  reg        [65:0]   _zz_io_input_payload_op1_10;
  reg        [65:0]   _zz_io_input_payload_op2_10;
  wire       [65:0]   _zz_io_input_payload_op1_11;
  wire       [65:0]   _zz_io_input_payload_op2_11;
  wire       [32:0]   _zz_io_input_payload_op1_12;
  wire       [32:0]   _zz_io_input_payload_op1_13;
  wire       [32:0]   _zz_io_input_payload_op2_12;
  wire       [32:0]   _zz_io_input_payload_op2_13;
  reg                 _zz_io_input_valid_2;
  reg        [32:0]   _zz_io_input_payload_op1_14;
  reg        [32:0]   _zz_io_input_payload_op1_15;
  reg        [32:0]   _zz_io_input_payload_op2_14;
  reg        [32:0]   _zz_io_input_payload_op2_15;
  reg        [33:0]   _zz_io_input_payload_op1_16;
  reg        [33:0]   _zz_io_input_payload_op2_16;
  reg                 _zz_output_valid;
  reg        [65:0]   _zz_output_payload_res;
  reg        [65:0]   _zz_output_payload_res_1;
  reg        [66:0]   _zz_output_payload_res_2;
  reg                 _zz_output_valid_1;
  reg        [131:0]  _zz_output_payload_res_3;
  wire       [65:0]   _zz_io_input_payload_op1_17;
  wire       [65:0]   _zz_io_input_payload_op2_17;
  wire       [32:0]   _zz_io_input_payload_op1_18;
  wire       [32:0]   _zz_io_input_payload_op1_19;
  wire       [32:0]   _zz_io_input_payload_op2_18;
  wire       [32:0]   _zz_io_input_payload_op2_19;
  reg                 _zz_io_input_valid_3;
  reg        [32:0]   _zz_io_input_payload_op1_20;
  reg        [32:0]   _zz_io_input_payload_op1_21;
  reg        [32:0]   _zz_io_input_payload_op2_20;
  reg        [32:0]   _zz_io_input_payload_op2_21;
  reg        [33:0]   _zz_io_input_payload_op1_22;
  reg        [33:0]   _zz_io_input_payload_op2_22;
  reg                 _zz_output_valid_2;
  reg        [65:0]   _zz_output_payload_res_4;
  reg        [65:0]   _zz_output_payload_res_5;
  reg        [66:0]   _zz_output_payload_res_6;
  reg                 _zz_output_valid_3;
  reg        [131:0]  _zz_output_payload_res_7;
  wire       [65:0]   _zz_io_input_payload_op1_23;
  wire       [65:0]   _zz_io_input_payload_op2_23;
  wire       [32:0]   _zz_io_input_payload_op1_24;
  wire       [32:0]   _zz_io_input_payload_op1_25;
  wire       [32:0]   _zz_io_input_payload_op2_24;
  wire       [32:0]   _zz_io_input_payload_op2_25;
  reg                 _zz_io_input_valid_4;
  reg        [32:0]   _zz_io_input_payload_op1_26;
  reg        [32:0]   _zz_io_input_payload_op1_27;
  reg        [32:0]   _zz_io_input_payload_op2_26;
  reg        [32:0]   _zz_io_input_payload_op2_27;
  reg        [33:0]   _zz_io_input_payload_op1_28;
  reg        [33:0]   _zz_io_input_payload_op2_28;
  reg                 _zz_output_valid_4;
  reg        [65:0]   _zz_output_payload_res_8;
  reg        [65:0]   _zz_output_payload_res_9;
  reg        [66:0]   _zz_output_payload_res_10;
  reg                 _zz_output_valid_5;
  reg        [131:0]  _zz_output_payload_res_11;
  reg                 _zz_output_valid_6;
  reg        [129:0]  _zz_output_payload_res_12;
  reg        [129:0]  _zz_output_payload_res_13;
  reg        [130:0]  _zz_output_payload_res_14;
  reg                 _zz_output_valid_7;
  reg        [257:0]  _zz_output_payload_res_15;
  wire       [128:0]  _zz_io_input_payload_op1_29;
  wire       [128:0]  _zz_io_input_payload_op2_29;
  wire       [64:0]   _zz_io_input_payload_op1_30;
  wire       [63:0]   _zz_io_input_payload_op1_31;
  wire       [64:0]   _zz_io_input_payload_op2_30;
  wire       [63:0]   _zz_io_input_payload_op2_31;
  reg                 _zz_io_input_valid_5;
  reg        [64:0]   _zz_io_input_payload_op1_32;
  reg        [63:0]   _zz_io_input_payload_op1_33;
  reg        [64:0]   _zz_io_input_payload_op2_32;
  reg        [63:0]   _zz_io_input_payload_op2_33;
  reg        [65:0]   _zz_io_input_payload_op1_34;
  reg        [65:0]   _zz_io_input_payload_op2_34;
  wire       [65:0]   _zz_io_input_payload_op1_35;
  wire       [65:0]   _zz_io_input_payload_op2_35;
  wire       [32:0]   _zz_io_input_payload_op1_36;
  wire       [32:0]   _zz_io_input_payload_op1_37;
  wire       [32:0]   _zz_io_input_payload_op2_36;
  wire       [32:0]   _zz_io_input_payload_op2_37;
  reg                 _zz_io_input_valid_6;
  reg        [32:0]   _zz_io_input_payload_op1_38;
  reg        [32:0]   _zz_io_input_payload_op1_39;
  reg        [32:0]   _zz_io_input_payload_op2_38;
  reg        [32:0]   _zz_io_input_payload_op2_39;
  reg        [33:0]   _zz_io_input_payload_op1_40;
  reg        [33:0]   _zz_io_input_payload_op2_40;
  reg                 _zz_output_valid_8;
  reg        [65:0]   _zz_output_payload_res_16;
  reg        [65:0]   _zz_output_payload_res_17;
  reg        [66:0]   _zz_output_payload_res_18;
  reg                 _zz_output_valid_9;
  reg        [131:0]  _zz_output_payload_res_19;
  wire       [65:0]   _zz_io_input_payload_op1_41;
  wire       [65:0]   _zz_io_input_payload_op2_41;
  wire       [32:0]   _zz_io_input_payload_op1_42;
  wire       [32:0]   _zz_io_input_payload_op1_43;
  wire       [32:0]   _zz_io_input_payload_op2_42;
  wire       [32:0]   _zz_io_input_payload_op2_43;
  reg                 _zz_io_input_valid_7;
  reg        [32:0]   _zz_io_input_payload_op1_44;
  reg        [32:0]   _zz_io_input_payload_op1_45;
  reg        [32:0]   _zz_io_input_payload_op2_44;
  reg        [32:0]   _zz_io_input_payload_op2_45;
  reg        [33:0]   _zz_io_input_payload_op1_46;
  reg        [33:0]   _zz_io_input_payload_op2_46;
  reg                 _zz_output_valid_10;
  reg        [65:0]   _zz_output_payload_res_20;
  reg        [65:0]   _zz_output_payload_res_21;
  reg        [66:0]   _zz_output_payload_res_22;
  reg                 _zz_output_valid_11;
  reg        [131:0]  _zz_output_payload_res_23;
  wire       [65:0]   _zz_io_input_payload_op1_47;
  wire       [65:0]   _zz_io_input_payload_op2_47;
  wire       [32:0]   _zz_io_input_payload_op1_48;
  wire       [32:0]   _zz_io_input_payload_op1_49;
  wire       [32:0]   _zz_io_input_payload_op2_48;
  wire       [32:0]   _zz_io_input_payload_op2_49;
  reg                 _zz_io_input_valid_8;
  reg        [32:0]   _zz_io_input_payload_op1_50;
  reg        [32:0]   _zz_io_input_payload_op1_51;
  reg        [32:0]   _zz_io_input_payload_op2_50;
  reg        [32:0]   _zz_io_input_payload_op2_51;
  reg        [33:0]   _zz_io_input_payload_op1_52;
  reg        [33:0]   _zz_io_input_payload_op2_52;
  reg                 _zz_output_valid_12;
  reg        [65:0]   _zz_output_payload_res_24;
  reg        [65:0]   _zz_output_payload_res_25;
  reg        [66:0]   _zz_output_payload_res_26;
  reg                 _zz_output_valid_13;
  reg        [131:0]  _zz_output_payload_res_27;
  reg                 _zz_output_valid_14;
  reg        [129:0]  _zz_output_payload_res_28;
  reg        [129:0]  _zz_output_payload_res_29;
  reg        [130:0]  _zz_output_payload_res_30;
  reg                 _zz_output_valid_15;
  reg        [257:0]  _zz_output_payload_res_31;
  wire       [128:0]  _zz_io_input_payload_op1_53;
  wire       [128:0]  _zz_io_input_payload_op2_53;
  wire       [64:0]   _zz_io_input_payload_op1_54;
  wire       [63:0]   _zz_io_input_payload_op1_55;
  wire       [64:0]   _zz_io_input_payload_op2_54;
  wire       [63:0]   _zz_io_input_payload_op2_55;
  reg                 _zz_io_input_valid_9;
  reg        [64:0]   _zz_io_input_payload_op1_56;
  reg        [63:0]   _zz_io_input_payload_op1_57;
  reg        [64:0]   _zz_io_input_payload_op2_56;
  reg        [63:0]   _zz_io_input_payload_op2_57;
  reg        [65:0]   _zz_io_input_payload_op1_58;
  reg        [65:0]   _zz_io_input_payload_op2_58;
  wire       [65:0]   _zz_io_input_payload_op1_59;
  wire       [65:0]   _zz_io_input_payload_op2_59;
  wire       [32:0]   _zz_io_input_payload_op1_60;
  wire       [32:0]   _zz_io_input_payload_op1_61;
  wire       [32:0]   _zz_io_input_payload_op2_60;
  wire       [32:0]   _zz_io_input_payload_op2_61;
  reg                 _zz_io_input_valid_10;
  reg        [32:0]   _zz_io_input_payload_op1_62;
  reg        [32:0]   _zz_io_input_payload_op1_63;
  reg        [32:0]   _zz_io_input_payload_op2_62;
  reg        [32:0]   _zz_io_input_payload_op2_63;
  reg        [33:0]   _zz_io_input_payload_op1_64;
  reg        [33:0]   _zz_io_input_payload_op2_64;
  reg                 _zz_output_valid_16;
  reg        [65:0]   _zz_output_payload_res_32;
  reg        [65:0]   _zz_output_payload_res_33;
  reg        [66:0]   _zz_output_payload_res_34;
  reg                 _zz_output_valid_17;
  reg        [131:0]  _zz_output_payload_res_35;
  wire       [65:0]   _zz_io_input_payload_op1_65;
  wire       [65:0]   _zz_io_input_payload_op2_65;
  wire       [32:0]   _zz_io_input_payload_op1_66;
  wire       [32:0]   _zz_io_input_payload_op1_67;
  wire       [32:0]   _zz_io_input_payload_op2_66;
  wire       [32:0]   _zz_io_input_payload_op2_67;
  reg                 _zz_io_input_valid_11;
  reg        [32:0]   _zz_io_input_payload_op1_68;
  reg        [32:0]   _zz_io_input_payload_op1_69;
  reg        [32:0]   _zz_io_input_payload_op2_68;
  reg        [32:0]   _zz_io_input_payload_op2_69;
  reg        [33:0]   _zz_io_input_payload_op1_70;
  reg        [33:0]   _zz_io_input_payload_op2_70;
  reg                 _zz_output_valid_18;
  reg        [65:0]   _zz_output_payload_res_36;
  reg        [65:0]   _zz_output_payload_res_37;
  reg        [66:0]   _zz_output_payload_res_38;
  reg                 _zz_output_valid_19;
  reg        [131:0]  _zz_output_payload_res_39;
  wire       [65:0]   _zz_io_input_payload_op1_71;
  wire       [65:0]   _zz_io_input_payload_op2_71;
  wire       [32:0]   _zz_io_input_payload_op1_72;
  wire       [32:0]   _zz_io_input_payload_op1_73;
  wire       [32:0]   _zz_io_input_payload_op2_72;
  wire       [32:0]   _zz_io_input_payload_op2_73;
  reg                 _zz_io_input_valid_12;
  reg        [32:0]   _zz_io_input_payload_op1_74;
  reg        [32:0]   _zz_io_input_payload_op1_75;
  reg        [32:0]   _zz_io_input_payload_op2_74;
  reg        [32:0]   _zz_io_input_payload_op2_75;
  reg        [33:0]   _zz_io_input_payload_op1_76;
  reg        [33:0]   _zz_io_input_payload_op2_76;
  reg                 _zz_output_valid_20;
  reg        [65:0]   _zz_output_payload_res_40;
  reg        [65:0]   _zz_output_payload_res_41;
  reg        [66:0]   _zz_output_payload_res_42;
  reg                 _zz_output_valid_21;
  reg        [131:0]  _zz_output_payload_res_43;
  reg                 _zz_output_valid_22;
  reg        [129:0]  _zz_output_payload_res_44;
  reg        [129:0]  _zz_output_payload_res_45;
  reg        [130:0]  _zz_output_payload_res_46;
  reg                 _zz_output_valid_23;
  reg        [257:0]  _zz_output_payload_res_47;
  reg                 _zz_output_valid_24;
  reg        [255:0]  _zz_output_payload_res_48;
  reg        [255:0]  _zz_output_payload_res_49;
  reg        [256:0]  _zz_output_payload_res_50;
  reg                 output_valid;
  reg        [511:0]  output_payload_res;

  assign _zz__zz_io_input_payload_op1_10_1 = {1'b0,_zz_io_input_payload_op1_7};
  assign _zz__zz_io_input_payload_op1_10 = {1'd0, _zz__zz_io_input_payload_op1_10_1};
  assign _zz__zz_io_input_payload_op2_10_1 = {1'b0,_zz_io_input_payload_op2_7};
  assign _zz__zz_io_input_payload_op2_10 = {1'd0, _zz__zz_io_input_payload_op2_10_1};
  assign _zz__zz_output_payload_res_2 = (_zz__zz_output_payload_res_2_1 - multiplierIPFlow_1216_io_output_payload_res);
  assign _zz__zz_output_payload_res_2_1 = (multiplierIPFlow_1217_io_output_payload_res - multiplierIPFlow_1215_io_output_payload_res);
  assign _zz__zz_output_payload_res_3 = (_zz__zz_output_payload_res_3_1 + _zz__zz_output_payload_res_3_2);
  assign _zz__zz_output_payload_res_3_1 = ({66'd0,_zz_output_payload_res} <<< 66);
  assign _zz__zz_output_payload_res_3_2 = {66'd0, _zz_output_payload_res_1};
  assign _zz__zz_output_payload_res_3_4 = ({33'd0,_zz_output_payload_res_2} <<< 33);
  assign _zz__zz_output_payload_res_3_3 = {32'd0, _zz__zz_output_payload_res_3_4};
  assign _zz__zz_output_payload_res_6 = (_zz__zz_output_payload_res_6_1 - multiplierIPFlow_1219_io_output_payload_res);
  assign _zz__zz_output_payload_res_6_1 = (multiplierIPFlow_1220_io_output_payload_res - multiplierIPFlow_1218_io_output_payload_res);
  assign _zz__zz_output_payload_res_7 = (_zz__zz_output_payload_res_7_1 + _zz__zz_output_payload_res_7_2);
  assign _zz__zz_output_payload_res_7_1 = ({66'd0,_zz_output_payload_res_4} <<< 66);
  assign _zz__zz_output_payload_res_7_2 = {66'd0, _zz_output_payload_res_5};
  assign _zz__zz_output_payload_res_7_4 = ({33'd0,_zz_output_payload_res_6} <<< 33);
  assign _zz__zz_output_payload_res_7_3 = {32'd0, _zz__zz_output_payload_res_7_4};
  assign _zz__zz_output_payload_res_10 = (_zz__zz_output_payload_res_10_1 - multiplierIPFlow_1222_io_output_payload_res);
  assign _zz__zz_output_payload_res_10_1 = (multiplierIPFlow_1223_io_output_payload_res - multiplierIPFlow_1221_io_output_payload_res);
  assign _zz__zz_output_payload_res_11 = (_zz__zz_output_payload_res_11_1 + _zz__zz_output_payload_res_11_2);
  assign _zz__zz_output_payload_res_11_1 = ({66'd0,_zz_output_payload_res_8} <<< 66);
  assign _zz__zz_output_payload_res_11_2 = {66'd0, _zz_output_payload_res_9};
  assign _zz__zz_output_payload_res_11_4 = ({33'd0,_zz_output_payload_res_10} <<< 33);
  assign _zz__zz_output_payload_res_11_3 = {32'd0, _zz__zz_output_payload_res_11_4};
  assign _zz__zz_output_payload_res_14 = (_zz__zz_output_payload_res_14_1 - _zz_output_payload_res_7);
  assign _zz__zz_output_payload_res_14_1 = (_zz_output_payload_res_11 - _zz_output_payload_res_3);
  assign _zz__zz_output_payload_res_15 = (_zz__zz_output_payload_res_15_1 + _zz__zz_output_payload_res_15_4);
  assign _zz__zz_output_payload_res_15_1 = (_zz__zz_output_payload_res_15_2 + _zz__zz_output_payload_res_15_3);
  assign _zz__zz_output_payload_res_15_2 = ({130'd0,_zz_output_payload_res_12} <<< 130);
  assign _zz__zz_output_payload_res_15_3 = {130'd0, _zz_output_payload_res_13};
  assign _zz__zz_output_payload_res_15_5 = ({65'd0,_zz_output_payload_res_14} <<< 65);
  assign _zz__zz_output_payload_res_15_4 = {64'd0, _zz__zz_output_payload_res_15_5};
  assign _zz__zz_io_input_payload_op1_34_1 = {1'b0,_zz_io_input_payload_op1_31};
  assign _zz__zz_io_input_payload_op1_34 = {1'd0, _zz__zz_io_input_payload_op1_34_1};
  assign _zz__zz_io_input_payload_op2_34_1 = {1'b0,_zz_io_input_payload_op2_31};
  assign _zz__zz_io_input_payload_op2_34 = {1'd0, _zz__zz_io_input_payload_op2_34_1};
  assign _zz__zz_output_payload_res_18 = (_zz__zz_output_payload_res_18_1 - multiplierIPFlow_1225_io_output_payload_res);
  assign _zz__zz_output_payload_res_18_1 = (multiplierIPFlow_1226_io_output_payload_res - multiplierIPFlow_1224_io_output_payload_res);
  assign _zz__zz_output_payload_res_19 = (_zz__zz_output_payload_res_19_1 + _zz__zz_output_payload_res_19_2);
  assign _zz__zz_output_payload_res_19_1 = ({66'd0,_zz_output_payload_res_16} <<< 66);
  assign _zz__zz_output_payload_res_19_2 = {66'd0, _zz_output_payload_res_17};
  assign _zz__zz_output_payload_res_19_4 = ({33'd0,_zz_output_payload_res_18} <<< 33);
  assign _zz__zz_output_payload_res_19_3 = {32'd0, _zz__zz_output_payload_res_19_4};
  assign _zz__zz_output_payload_res_22 = (_zz__zz_output_payload_res_22_1 - multiplierIPFlow_1228_io_output_payload_res);
  assign _zz__zz_output_payload_res_22_1 = (multiplierIPFlow_1229_io_output_payload_res - multiplierIPFlow_1227_io_output_payload_res);
  assign _zz__zz_output_payload_res_23 = (_zz__zz_output_payload_res_23_1 + _zz__zz_output_payload_res_23_2);
  assign _zz__zz_output_payload_res_23_1 = ({66'd0,_zz_output_payload_res_20} <<< 66);
  assign _zz__zz_output_payload_res_23_2 = {66'd0, _zz_output_payload_res_21};
  assign _zz__zz_output_payload_res_23_4 = ({33'd0,_zz_output_payload_res_22} <<< 33);
  assign _zz__zz_output_payload_res_23_3 = {32'd0, _zz__zz_output_payload_res_23_4};
  assign _zz__zz_output_payload_res_26 = (_zz__zz_output_payload_res_26_1 - multiplierIPFlow_1231_io_output_payload_res);
  assign _zz__zz_output_payload_res_26_1 = (multiplierIPFlow_1232_io_output_payload_res - multiplierIPFlow_1230_io_output_payload_res);
  assign _zz__zz_output_payload_res_27 = (_zz__zz_output_payload_res_27_1 + _zz__zz_output_payload_res_27_2);
  assign _zz__zz_output_payload_res_27_1 = ({66'd0,_zz_output_payload_res_24} <<< 66);
  assign _zz__zz_output_payload_res_27_2 = {66'd0, _zz_output_payload_res_25};
  assign _zz__zz_output_payload_res_27_4 = ({33'd0,_zz_output_payload_res_26} <<< 33);
  assign _zz__zz_output_payload_res_27_3 = {32'd0, _zz__zz_output_payload_res_27_4};
  assign _zz__zz_output_payload_res_30 = (_zz__zz_output_payload_res_30_1 - _zz_output_payload_res_23);
  assign _zz__zz_output_payload_res_30_1 = (_zz_output_payload_res_27 - _zz_output_payload_res_19);
  assign _zz__zz_output_payload_res_31 = (_zz__zz_output_payload_res_31_1 + _zz__zz_output_payload_res_31_4);
  assign _zz__zz_output_payload_res_31_1 = (_zz__zz_output_payload_res_31_2 + _zz__zz_output_payload_res_31_3);
  assign _zz__zz_output_payload_res_31_2 = ({130'd0,_zz_output_payload_res_28} <<< 130);
  assign _zz__zz_output_payload_res_31_3 = {130'd0, _zz_output_payload_res_29};
  assign _zz__zz_output_payload_res_31_5 = ({65'd0,_zz_output_payload_res_30} <<< 65);
  assign _zz__zz_output_payload_res_31_4 = {64'd0, _zz__zz_output_payload_res_31_5};
  assign _zz__zz_io_input_payload_op1_58_1 = {1'b0,_zz_io_input_payload_op1_55};
  assign _zz__zz_io_input_payload_op1_58 = {1'd0, _zz__zz_io_input_payload_op1_58_1};
  assign _zz__zz_io_input_payload_op2_58_1 = {1'b0,_zz_io_input_payload_op2_55};
  assign _zz__zz_io_input_payload_op2_58 = {1'd0, _zz__zz_io_input_payload_op2_58_1};
  assign _zz__zz_output_payload_res_34 = (_zz__zz_output_payload_res_34_1 - multiplierIPFlow_1234_io_output_payload_res);
  assign _zz__zz_output_payload_res_34_1 = (multiplierIPFlow_1235_io_output_payload_res - multiplierIPFlow_1233_io_output_payload_res);
  assign _zz__zz_output_payload_res_35 = (_zz__zz_output_payload_res_35_1 + _zz__zz_output_payload_res_35_2);
  assign _zz__zz_output_payload_res_35_1 = ({66'd0,_zz_output_payload_res_32} <<< 66);
  assign _zz__zz_output_payload_res_35_2 = {66'd0, _zz_output_payload_res_33};
  assign _zz__zz_output_payload_res_35_4 = ({33'd0,_zz_output_payload_res_34} <<< 33);
  assign _zz__zz_output_payload_res_35_3 = {32'd0, _zz__zz_output_payload_res_35_4};
  assign _zz__zz_output_payload_res_38 = (_zz__zz_output_payload_res_38_1 - multiplierIPFlow_1237_io_output_payload_res);
  assign _zz__zz_output_payload_res_38_1 = (multiplierIPFlow_1238_io_output_payload_res - multiplierIPFlow_1236_io_output_payload_res);
  assign _zz__zz_output_payload_res_39 = (_zz__zz_output_payload_res_39_1 + _zz__zz_output_payload_res_39_2);
  assign _zz__zz_output_payload_res_39_1 = ({66'd0,_zz_output_payload_res_36} <<< 66);
  assign _zz__zz_output_payload_res_39_2 = {66'd0, _zz_output_payload_res_37};
  assign _zz__zz_output_payload_res_39_4 = ({33'd0,_zz_output_payload_res_38} <<< 33);
  assign _zz__zz_output_payload_res_39_3 = {32'd0, _zz__zz_output_payload_res_39_4};
  assign _zz__zz_output_payload_res_42 = (_zz__zz_output_payload_res_42_1 - multiplierIPFlow_1240_io_output_payload_res);
  assign _zz__zz_output_payload_res_42_1 = (multiplierIPFlow_1241_io_output_payload_res - multiplierIPFlow_1239_io_output_payload_res);
  assign _zz__zz_output_payload_res_43 = (_zz__zz_output_payload_res_43_1 + _zz__zz_output_payload_res_43_2);
  assign _zz__zz_output_payload_res_43_1 = ({66'd0,_zz_output_payload_res_40} <<< 66);
  assign _zz__zz_output_payload_res_43_2 = {66'd0, _zz_output_payload_res_41};
  assign _zz__zz_output_payload_res_43_4 = ({33'd0,_zz_output_payload_res_42} <<< 33);
  assign _zz__zz_output_payload_res_43_3 = {32'd0, _zz__zz_output_payload_res_43_4};
  assign _zz__zz_output_payload_res_46 = (_zz__zz_output_payload_res_46_1 - _zz_output_payload_res_39);
  assign _zz__zz_output_payload_res_46_1 = (_zz_output_payload_res_43 - _zz_output_payload_res_35);
  assign _zz__zz_output_payload_res_47 = (_zz__zz_output_payload_res_47_1 + _zz__zz_output_payload_res_47_4);
  assign _zz__zz_output_payload_res_47_1 = (_zz__zz_output_payload_res_47_2 + _zz__zz_output_payload_res_47_3);
  assign _zz__zz_output_payload_res_47_2 = ({130'd0,_zz_output_payload_res_44} <<< 130);
  assign _zz__zz_output_payload_res_47_3 = {130'd0, _zz_output_payload_res_45};
  assign _zz__zz_output_payload_res_47_5 = ({65'd0,_zz_output_payload_res_46} <<< 65);
  assign _zz__zz_output_payload_res_47_4 = {64'd0, _zz__zz_output_payload_res_47_5};
  assign _zz__zz_output_payload_res_50 = (_zz__zz_output_payload_res_50_1 - _zz_output_payload_res_31);
  assign _zz__zz_output_payload_res_50_1 = (_zz_output_payload_res_47 - _zz_output_payload_res_15);
  assign _zz_output_payload_res_51 = (_zz_output_payload_res_52 + _zz_output_payload_res_53);
  assign _zz_output_payload_res_52 = ({256'd0,_zz_output_payload_res_48} <<< 256);
  assign _zz_output_payload_res_53 = {256'd0, _zz_output_payload_res_49};
  assign _zz_output_payload_res_55 = ({128'd0,_zz_output_payload_res_50} <<< 128);
  assign _zz_output_payload_res_54 = {127'd0, _zz_output_payload_res_55};
  MultiplierIPFlow multiplierIPFlow_1215 (
    .io_input_valid           (_zz_io_input_valid_2                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1215_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1215_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1215_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1215_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1216 (
    .io_input_valid           (_zz_io_input_valid_2                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1216_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1216_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1216_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1216_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1217 (
    .io_input_valid           (_zz_io_input_valid_2                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_16[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_16[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1217_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1217_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1218 (
    .io_input_valid           (_zz_io_input_valid_3                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1218_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1218_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1218_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1218_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1219 (
    .io_input_valid           (_zz_io_input_valid_3                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1219_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1219_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1219_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1219_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1220 (
    .io_input_valid           (_zz_io_input_valid_3                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_22[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_22[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1220_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1220_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1221 (
    .io_input_valid           (_zz_io_input_valid_4                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1221_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1221_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1221_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1221_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1222 (
    .io_input_valid           (_zz_io_input_valid_4                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1222_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1222_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1222_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1222_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1223 (
    .io_input_valid           (_zz_io_input_valid_4                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_28[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_28[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1223_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1223_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1224 (
    .io_input_valid           (_zz_io_input_valid_6                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1224_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1224_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1224_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1224_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1225 (
    .io_input_valid           (_zz_io_input_valid_6                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1225_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1225_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1225_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1225_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1226 (
    .io_input_valid           (_zz_io_input_valid_6                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_40[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_40[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1226_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1226_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1227 (
    .io_input_valid           (_zz_io_input_valid_7                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1227_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1227_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1227_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1227_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1228 (
    .io_input_valid           (_zz_io_input_valid_7                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1228_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1228_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1228_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1228_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1229 (
    .io_input_valid           (_zz_io_input_valid_7                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_46[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_46[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1229_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1229_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1230 (
    .io_input_valid           (_zz_io_input_valid_8                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1230_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1230_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1230_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1230_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1231 (
    .io_input_valid           (_zz_io_input_valid_8                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1231_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1231_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1231_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1231_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1232 (
    .io_input_valid           (_zz_io_input_valid_8                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_52[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_52[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1232_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1232_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1233 (
    .io_input_valid           (_zz_io_input_valid_10                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1233_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1233_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1233_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1233_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1234 (
    .io_input_valid           (_zz_io_input_valid_10                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1234_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1234_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1234_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1234_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1235 (
    .io_input_valid           (_zz_io_input_valid_10                              ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_64[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_64[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1235_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1235_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1236 (
    .io_input_valid           (_zz_io_input_valid_11                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1236_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1236_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1236_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1236_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1237 (
    .io_input_valid           (_zz_io_input_valid_11                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1237_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1237_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1237_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1237_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1238 (
    .io_input_valid           (_zz_io_input_valid_11                              ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_70[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_70[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1238_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1238_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1239 (
    .io_input_valid           (_zz_io_input_valid_12                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1239_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1239_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1239_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1239_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1240 (
    .io_input_valid           (_zz_io_input_valid_12                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1240_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1240_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1240_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1240_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1241 (
    .io_input_valid           (_zz_io_input_valid_12                              ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_76[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_76[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1241_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1241_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  assign _zz_io_input_payload_op1 = io_input_payload_op1[127 : 0];
  assign _zz_io_input_payload_op1_1 = io_input_payload_op1[255 : 128];
  assign _zz_io_input_payload_op2 = io_input_payload_op2[127 : 0];
  assign _zz_io_input_payload_op2_1 = io_input_payload_op2[255 : 128];
  assign _zz_io_input_payload_op1_5 = {1'd0, _zz_io_input_payload_op1_3};
  assign _zz_io_input_payload_op2_5 = {1'd0, _zz_io_input_payload_op2_3};
  assign _zz_io_input_payload_op1_6 = _zz_io_input_payload_op1_5[64 : 0];
  assign _zz_io_input_payload_op1_7 = _zz_io_input_payload_op1_5[128 : 65];
  assign _zz_io_input_payload_op2_6 = _zz_io_input_payload_op2_5[64 : 0];
  assign _zz_io_input_payload_op2_7 = _zz_io_input_payload_op2_5[128 : 65];
  assign _zz_io_input_payload_op1_11 = {2'd0, _zz_io_input_payload_op1_9};
  assign _zz_io_input_payload_op2_11 = {2'd0, _zz_io_input_payload_op2_9};
  assign _zz_io_input_payload_op1_12 = _zz_io_input_payload_op1_11[32 : 0];
  assign _zz_io_input_payload_op1_13 = _zz_io_input_payload_op1_11[65 : 33];
  assign _zz_io_input_payload_op2_12 = _zz_io_input_payload_op2_11[32 : 0];
  assign _zz_io_input_payload_op2_13 = _zz_io_input_payload_op2_11[65 : 33];
  assign multiplierIPFlow_1215_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_15};
  assign multiplierIPFlow_1215_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_15};
  assign multiplierIPFlow_1216_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_14};
  assign multiplierIPFlow_1216_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_14};
  assign _zz_io_input_payload_op1_17 = {1'd0, _zz_io_input_payload_op1_8};
  assign _zz_io_input_payload_op2_17 = {1'd0, _zz_io_input_payload_op2_8};
  assign _zz_io_input_payload_op1_18 = _zz_io_input_payload_op1_17[32 : 0];
  assign _zz_io_input_payload_op1_19 = _zz_io_input_payload_op1_17[65 : 33];
  assign _zz_io_input_payload_op2_18 = _zz_io_input_payload_op2_17[32 : 0];
  assign _zz_io_input_payload_op2_19 = _zz_io_input_payload_op2_17[65 : 33];
  assign multiplierIPFlow_1218_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_21};
  assign multiplierIPFlow_1218_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_21};
  assign multiplierIPFlow_1219_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_20};
  assign multiplierIPFlow_1219_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_20};
  assign _zz_io_input_payload_op1_23 = _zz_io_input_payload_op1_10;
  assign _zz_io_input_payload_op2_23 = _zz_io_input_payload_op2_10;
  assign _zz_io_input_payload_op1_24 = _zz_io_input_payload_op1_23[32 : 0];
  assign _zz_io_input_payload_op1_25 = _zz_io_input_payload_op1_23[65 : 33];
  assign _zz_io_input_payload_op2_24 = _zz_io_input_payload_op2_23[32 : 0];
  assign _zz_io_input_payload_op2_25 = _zz_io_input_payload_op2_23[65 : 33];
  assign multiplierIPFlow_1221_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_27};
  assign multiplierIPFlow_1221_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_27};
  assign multiplierIPFlow_1222_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_26};
  assign multiplierIPFlow_1222_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_26};
  assign _zz_io_input_payload_op1_29 = {1'd0, _zz_io_input_payload_op1_2};
  assign _zz_io_input_payload_op2_29 = {1'd0, _zz_io_input_payload_op2_2};
  assign _zz_io_input_payload_op1_30 = _zz_io_input_payload_op1_29[64 : 0];
  assign _zz_io_input_payload_op1_31 = _zz_io_input_payload_op1_29[128 : 65];
  assign _zz_io_input_payload_op2_30 = _zz_io_input_payload_op2_29[64 : 0];
  assign _zz_io_input_payload_op2_31 = _zz_io_input_payload_op2_29[128 : 65];
  assign _zz_io_input_payload_op1_35 = {2'd0, _zz_io_input_payload_op1_33};
  assign _zz_io_input_payload_op2_35 = {2'd0, _zz_io_input_payload_op2_33};
  assign _zz_io_input_payload_op1_36 = _zz_io_input_payload_op1_35[32 : 0];
  assign _zz_io_input_payload_op1_37 = _zz_io_input_payload_op1_35[65 : 33];
  assign _zz_io_input_payload_op2_36 = _zz_io_input_payload_op2_35[32 : 0];
  assign _zz_io_input_payload_op2_37 = _zz_io_input_payload_op2_35[65 : 33];
  assign multiplierIPFlow_1224_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_39};
  assign multiplierIPFlow_1224_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_39};
  assign multiplierIPFlow_1225_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_38};
  assign multiplierIPFlow_1225_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_38};
  assign _zz_io_input_payload_op1_41 = {1'd0, _zz_io_input_payload_op1_32};
  assign _zz_io_input_payload_op2_41 = {1'd0, _zz_io_input_payload_op2_32};
  assign _zz_io_input_payload_op1_42 = _zz_io_input_payload_op1_41[32 : 0];
  assign _zz_io_input_payload_op1_43 = _zz_io_input_payload_op1_41[65 : 33];
  assign _zz_io_input_payload_op2_42 = _zz_io_input_payload_op2_41[32 : 0];
  assign _zz_io_input_payload_op2_43 = _zz_io_input_payload_op2_41[65 : 33];
  assign multiplierIPFlow_1227_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_45};
  assign multiplierIPFlow_1227_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_45};
  assign multiplierIPFlow_1228_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_44};
  assign multiplierIPFlow_1228_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_44};
  assign _zz_io_input_payload_op1_47 = _zz_io_input_payload_op1_34;
  assign _zz_io_input_payload_op2_47 = _zz_io_input_payload_op2_34;
  assign _zz_io_input_payload_op1_48 = _zz_io_input_payload_op1_47[32 : 0];
  assign _zz_io_input_payload_op1_49 = _zz_io_input_payload_op1_47[65 : 33];
  assign _zz_io_input_payload_op2_48 = _zz_io_input_payload_op2_47[32 : 0];
  assign _zz_io_input_payload_op2_49 = _zz_io_input_payload_op2_47[65 : 33];
  assign multiplierIPFlow_1230_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_51};
  assign multiplierIPFlow_1230_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_51};
  assign multiplierIPFlow_1231_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_50};
  assign multiplierIPFlow_1231_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_50};
  assign _zz_io_input_payload_op1_53 = _zz_io_input_payload_op1_4;
  assign _zz_io_input_payload_op2_53 = _zz_io_input_payload_op2_4;
  assign _zz_io_input_payload_op1_54 = _zz_io_input_payload_op1_53[64 : 0];
  assign _zz_io_input_payload_op1_55 = _zz_io_input_payload_op1_53[128 : 65];
  assign _zz_io_input_payload_op2_54 = _zz_io_input_payload_op2_53[64 : 0];
  assign _zz_io_input_payload_op2_55 = _zz_io_input_payload_op2_53[128 : 65];
  assign _zz_io_input_payload_op1_59 = {2'd0, _zz_io_input_payload_op1_57};
  assign _zz_io_input_payload_op2_59 = {2'd0, _zz_io_input_payload_op2_57};
  assign _zz_io_input_payload_op1_60 = _zz_io_input_payload_op1_59[32 : 0];
  assign _zz_io_input_payload_op1_61 = _zz_io_input_payload_op1_59[65 : 33];
  assign _zz_io_input_payload_op2_60 = _zz_io_input_payload_op2_59[32 : 0];
  assign _zz_io_input_payload_op2_61 = _zz_io_input_payload_op2_59[65 : 33];
  assign multiplierIPFlow_1233_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_63};
  assign multiplierIPFlow_1233_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_63};
  assign multiplierIPFlow_1234_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_62};
  assign multiplierIPFlow_1234_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_62};
  assign _zz_io_input_payload_op1_65 = {1'd0, _zz_io_input_payload_op1_56};
  assign _zz_io_input_payload_op2_65 = {1'd0, _zz_io_input_payload_op2_56};
  assign _zz_io_input_payload_op1_66 = _zz_io_input_payload_op1_65[32 : 0];
  assign _zz_io_input_payload_op1_67 = _zz_io_input_payload_op1_65[65 : 33];
  assign _zz_io_input_payload_op2_66 = _zz_io_input_payload_op2_65[32 : 0];
  assign _zz_io_input_payload_op2_67 = _zz_io_input_payload_op2_65[65 : 33];
  assign multiplierIPFlow_1236_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_69};
  assign multiplierIPFlow_1236_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_69};
  assign multiplierIPFlow_1237_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_68};
  assign multiplierIPFlow_1237_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_68};
  assign _zz_io_input_payload_op1_71 = _zz_io_input_payload_op1_58;
  assign _zz_io_input_payload_op2_71 = _zz_io_input_payload_op2_58;
  assign _zz_io_input_payload_op1_72 = _zz_io_input_payload_op1_71[32 : 0];
  assign _zz_io_input_payload_op1_73 = _zz_io_input_payload_op1_71[65 : 33];
  assign _zz_io_input_payload_op2_72 = _zz_io_input_payload_op2_71[32 : 0];
  assign _zz_io_input_payload_op2_73 = _zz_io_input_payload_op2_71[65 : 33];
  assign multiplierIPFlow_1239_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_75};
  assign multiplierIPFlow_1239_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_75};
  assign multiplierIPFlow_1240_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_74};
  assign multiplierIPFlow_1240_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_74};
  assign io_output_valid = output_valid;
  assign io_output_payload_res = output_payload_res;
  always @(posedge clk) begin
    if(!resetn) begin
      _zz_io_input_valid <= 1'b0;
      _zz_io_input_valid_1 <= 1'b0;
      _zz_io_input_valid_2 <= 1'b0;
      _zz_output_valid <= 1'b0;
      _zz_output_valid_1 <= 1'b0;
      _zz_io_input_valid_3 <= 1'b0;
      _zz_output_valid_2 <= 1'b0;
      _zz_output_valid_3 <= 1'b0;
      _zz_io_input_valid_4 <= 1'b0;
      _zz_output_valid_4 <= 1'b0;
      _zz_output_valid_5 <= 1'b0;
      _zz_output_valid_6 <= 1'b0;
      _zz_output_valid_7 <= 1'b0;
      _zz_io_input_valid_5 <= 1'b0;
      _zz_io_input_valid_6 <= 1'b0;
      _zz_output_valid_8 <= 1'b0;
      _zz_output_valid_9 <= 1'b0;
      _zz_io_input_valid_7 <= 1'b0;
      _zz_output_valid_10 <= 1'b0;
      _zz_output_valid_11 <= 1'b0;
      _zz_io_input_valid_8 <= 1'b0;
      _zz_output_valid_12 <= 1'b0;
      _zz_output_valid_13 <= 1'b0;
      _zz_output_valid_14 <= 1'b0;
      _zz_output_valid_15 <= 1'b0;
      _zz_io_input_valid_9 <= 1'b0;
      _zz_io_input_valid_10 <= 1'b0;
      _zz_output_valid_16 <= 1'b0;
      _zz_output_valid_17 <= 1'b0;
      _zz_io_input_valid_11 <= 1'b0;
      _zz_output_valid_18 <= 1'b0;
      _zz_output_valid_19 <= 1'b0;
      _zz_io_input_valid_12 <= 1'b0;
      _zz_output_valid_20 <= 1'b0;
      _zz_output_valid_21 <= 1'b0;
      _zz_output_valid_22 <= 1'b0;
      _zz_output_valid_23 <= 1'b0;
      _zz_output_valid_24 <= 1'b0;
      output_valid <= 1'b0;
    end else begin
      _zz_io_input_valid <= io_input_valid;
      _zz_io_input_valid_1 <= _zz_io_input_valid;
      _zz_io_input_valid_2 <= _zz_io_input_valid_1;
      _zz_output_valid <= ((multiplierIPFlow_1215_io_output_valid && multiplierIPFlow_1216_io_output_valid) && multiplierIPFlow_1217_io_output_valid);
      _zz_output_valid_1 <= _zz_output_valid;
      _zz_io_input_valid_3 <= _zz_io_input_valid_1;
      _zz_output_valid_2 <= ((multiplierIPFlow_1218_io_output_valid && multiplierIPFlow_1219_io_output_valid) && multiplierIPFlow_1220_io_output_valid);
      _zz_output_valid_3 <= _zz_output_valid_2;
      _zz_io_input_valid_4 <= _zz_io_input_valid_1;
      _zz_output_valid_4 <= ((multiplierIPFlow_1221_io_output_valid && multiplierIPFlow_1222_io_output_valid) && multiplierIPFlow_1223_io_output_valid);
      _zz_output_valid_5 <= _zz_output_valid_4;
      _zz_output_valid_6 <= ((_zz_output_valid_1 && _zz_output_valid_3) && _zz_output_valid_5);
      _zz_output_valid_7 <= _zz_output_valid_6;
      _zz_io_input_valid_5 <= _zz_io_input_valid;
      _zz_io_input_valid_6 <= _zz_io_input_valid_5;
      _zz_output_valid_8 <= ((multiplierIPFlow_1224_io_output_valid && multiplierIPFlow_1225_io_output_valid) && multiplierIPFlow_1226_io_output_valid);
      _zz_output_valid_9 <= _zz_output_valid_8;
      _zz_io_input_valid_7 <= _zz_io_input_valid_5;
      _zz_output_valid_10 <= ((multiplierIPFlow_1227_io_output_valid && multiplierIPFlow_1228_io_output_valid) && multiplierIPFlow_1229_io_output_valid);
      _zz_output_valid_11 <= _zz_output_valid_10;
      _zz_io_input_valid_8 <= _zz_io_input_valid_5;
      _zz_output_valid_12 <= ((multiplierIPFlow_1230_io_output_valid && multiplierIPFlow_1231_io_output_valid) && multiplierIPFlow_1232_io_output_valid);
      _zz_output_valid_13 <= _zz_output_valid_12;
      _zz_output_valid_14 <= ((_zz_output_valid_9 && _zz_output_valid_11) && _zz_output_valid_13);
      _zz_output_valid_15 <= _zz_output_valid_14;
      _zz_io_input_valid_9 <= _zz_io_input_valid;
      _zz_io_input_valid_10 <= _zz_io_input_valid_9;
      _zz_output_valid_16 <= ((multiplierIPFlow_1233_io_output_valid && multiplierIPFlow_1234_io_output_valid) && multiplierIPFlow_1235_io_output_valid);
      _zz_output_valid_17 <= _zz_output_valid_16;
      _zz_io_input_valid_11 <= _zz_io_input_valid_9;
      _zz_output_valid_18 <= ((multiplierIPFlow_1236_io_output_valid && multiplierIPFlow_1237_io_output_valid) && multiplierIPFlow_1238_io_output_valid);
      _zz_output_valid_19 <= _zz_output_valid_18;
      _zz_io_input_valid_12 <= _zz_io_input_valid_9;
      _zz_output_valid_20 <= ((multiplierIPFlow_1239_io_output_valid && multiplierIPFlow_1240_io_output_valid) && multiplierIPFlow_1241_io_output_valid);
      _zz_output_valid_21 <= _zz_output_valid_20;
      _zz_output_valid_22 <= ((_zz_output_valid_17 && _zz_output_valid_19) && _zz_output_valid_21);
      _zz_output_valid_23 <= _zz_output_valid_22;
      _zz_output_valid_24 <= ((_zz_output_valid_7 && _zz_output_valid_15) && _zz_output_valid_23);
      output_valid <= _zz_output_valid_24;
    end
  end

  always @(posedge clk) begin
    _zz_io_input_payload_op1_2 <= _zz_io_input_payload_op1;
    _zz_io_input_payload_op1_3 <= _zz_io_input_payload_op1_1;
    _zz_io_input_payload_op2_2 <= _zz_io_input_payload_op2;
    _zz_io_input_payload_op2_3 <= _zz_io_input_payload_op2_1;
    _zz_io_input_payload_op1_4 <= ({1'b0,_zz_io_input_payload_op1} + {1'b0,_zz_io_input_payload_op1_1});
    _zz_io_input_payload_op2_4 <= ({1'b0,_zz_io_input_payload_op2} + {1'b0,_zz_io_input_payload_op2_1});
    _zz_io_input_payload_op1_8 <= _zz_io_input_payload_op1_6;
    _zz_io_input_payload_op1_9 <= _zz_io_input_payload_op1_7;
    _zz_io_input_payload_op2_8 <= _zz_io_input_payload_op2_6;
    _zz_io_input_payload_op2_9 <= _zz_io_input_payload_op2_7;
    _zz_io_input_payload_op1_10 <= ({1'b0,_zz_io_input_payload_op1_6} + _zz__zz_io_input_payload_op1_10);
    _zz_io_input_payload_op2_10 <= ({1'b0,_zz_io_input_payload_op2_6} + _zz__zz_io_input_payload_op2_10);
    _zz_io_input_payload_op1_14 <= _zz_io_input_payload_op1_12;
    _zz_io_input_payload_op1_15 <= _zz_io_input_payload_op1_13;
    _zz_io_input_payload_op2_14 <= _zz_io_input_payload_op2_12;
    _zz_io_input_payload_op2_15 <= _zz_io_input_payload_op2_13;
    _zz_io_input_payload_op1_16 <= ({1'b0,_zz_io_input_payload_op1_12} + {1'b0,_zz_io_input_payload_op1_13});
    _zz_io_input_payload_op2_16 <= ({1'b0,_zz_io_input_payload_op2_12} + {1'b0,_zz_io_input_payload_op2_13});
    _zz_output_payload_res <= multiplierIPFlow_1215_io_output_payload_res[65:0];
    _zz_output_payload_res_1 <= multiplierIPFlow_1216_io_output_payload_res[65:0];
    _zz_output_payload_res_2 <= _zz__zz_output_payload_res_2[66:0];
    _zz_output_payload_res_3 <= (_zz__zz_output_payload_res_3 + _zz__zz_output_payload_res_3_3);
    _zz_io_input_payload_op1_20 <= _zz_io_input_payload_op1_18;
    _zz_io_input_payload_op1_21 <= _zz_io_input_payload_op1_19;
    _zz_io_input_payload_op2_20 <= _zz_io_input_payload_op2_18;
    _zz_io_input_payload_op2_21 <= _zz_io_input_payload_op2_19;
    _zz_io_input_payload_op1_22 <= ({1'b0,_zz_io_input_payload_op1_18} + {1'b0,_zz_io_input_payload_op1_19});
    _zz_io_input_payload_op2_22 <= ({1'b0,_zz_io_input_payload_op2_18} + {1'b0,_zz_io_input_payload_op2_19});
    _zz_output_payload_res_4 <= multiplierIPFlow_1218_io_output_payload_res[65:0];
    _zz_output_payload_res_5 <= multiplierIPFlow_1219_io_output_payload_res[65:0];
    _zz_output_payload_res_6 <= _zz__zz_output_payload_res_6[66:0];
    _zz_output_payload_res_7 <= (_zz__zz_output_payload_res_7 + _zz__zz_output_payload_res_7_3);
    _zz_io_input_payload_op1_26 <= _zz_io_input_payload_op1_24;
    _zz_io_input_payload_op1_27 <= _zz_io_input_payload_op1_25;
    _zz_io_input_payload_op2_26 <= _zz_io_input_payload_op2_24;
    _zz_io_input_payload_op2_27 <= _zz_io_input_payload_op2_25;
    _zz_io_input_payload_op1_28 <= ({1'b0,_zz_io_input_payload_op1_24} + {1'b0,_zz_io_input_payload_op1_25});
    _zz_io_input_payload_op2_28 <= ({1'b0,_zz_io_input_payload_op2_24} + {1'b0,_zz_io_input_payload_op2_25});
    _zz_output_payload_res_8 <= multiplierIPFlow_1221_io_output_payload_res[65:0];
    _zz_output_payload_res_9 <= multiplierIPFlow_1222_io_output_payload_res[65:0];
    _zz_output_payload_res_10 <= _zz__zz_output_payload_res_10[66:0];
    _zz_output_payload_res_11 <= (_zz__zz_output_payload_res_11 + _zz__zz_output_payload_res_11_3);
    _zz_output_payload_res_12 <= _zz_output_payload_res_3[129:0];
    _zz_output_payload_res_13 <= _zz_output_payload_res_7[129:0];
    _zz_output_payload_res_14 <= _zz__zz_output_payload_res_14[130:0];
    _zz_output_payload_res_15 <= _zz__zz_output_payload_res_15[257:0];
    _zz_io_input_payload_op1_32 <= _zz_io_input_payload_op1_30;
    _zz_io_input_payload_op1_33 <= _zz_io_input_payload_op1_31;
    _zz_io_input_payload_op2_32 <= _zz_io_input_payload_op2_30;
    _zz_io_input_payload_op2_33 <= _zz_io_input_payload_op2_31;
    _zz_io_input_payload_op1_34 <= ({1'b0,_zz_io_input_payload_op1_30} + _zz__zz_io_input_payload_op1_34);
    _zz_io_input_payload_op2_34 <= ({1'b0,_zz_io_input_payload_op2_30} + _zz__zz_io_input_payload_op2_34);
    _zz_io_input_payload_op1_38 <= _zz_io_input_payload_op1_36;
    _zz_io_input_payload_op1_39 <= _zz_io_input_payload_op1_37;
    _zz_io_input_payload_op2_38 <= _zz_io_input_payload_op2_36;
    _zz_io_input_payload_op2_39 <= _zz_io_input_payload_op2_37;
    _zz_io_input_payload_op1_40 <= ({1'b0,_zz_io_input_payload_op1_36} + {1'b0,_zz_io_input_payload_op1_37});
    _zz_io_input_payload_op2_40 <= ({1'b0,_zz_io_input_payload_op2_36} + {1'b0,_zz_io_input_payload_op2_37});
    _zz_output_payload_res_16 <= multiplierIPFlow_1224_io_output_payload_res[65:0];
    _zz_output_payload_res_17 <= multiplierIPFlow_1225_io_output_payload_res[65:0];
    _zz_output_payload_res_18 <= _zz__zz_output_payload_res_18[66:0];
    _zz_output_payload_res_19 <= (_zz__zz_output_payload_res_19 + _zz__zz_output_payload_res_19_3);
    _zz_io_input_payload_op1_44 <= _zz_io_input_payload_op1_42;
    _zz_io_input_payload_op1_45 <= _zz_io_input_payload_op1_43;
    _zz_io_input_payload_op2_44 <= _zz_io_input_payload_op2_42;
    _zz_io_input_payload_op2_45 <= _zz_io_input_payload_op2_43;
    _zz_io_input_payload_op1_46 <= ({1'b0,_zz_io_input_payload_op1_42} + {1'b0,_zz_io_input_payload_op1_43});
    _zz_io_input_payload_op2_46 <= ({1'b0,_zz_io_input_payload_op2_42} + {1'b0,_zz_io_input_payload_op2_43});
    _zz_output_payload_res_20 <= multiplierIPFlow_1227_io_output_payload_res[65:0];
    _zz_output_payload_res_21 <= multiplierIPFlow_1228_io_output_payload_res[65:0];
    _zz_output_payload_res_22 <= _zz__zz_output_payload_res_22[66:0];
    _zz_output_payload_res_23 <= (_zz__zz_output_payload_res_23 + _zz__zz_output_payload_res_23_3);
    _zz_io_input_payload_op1_50 <= _zz_io_input_payload_op1_48;
    _zz_io_input_payload_op1_51 <= _zz_io_input_payload_op1_49;
    _zz_io_input_payload_op2_50 <= _zz_io_input_payload_op2_48;
    _zz_io_input_payload_op2_51 <= _zz_io_input_payload_op2_49;
    _zz_io_input_payload_op1_52 <= ({1'b0,_zz_io_input_payload_op1_48} + {1'b0,_zz_io_input_payload_op1_49});
    _zz_io_input_payload_op2_52 <= ({1'b0,_zz_io_input_payload_op2_48} + {1'b0,_zz_io_input_payload_op2_49});
    _zz_output_payload_res_24 <= multiplierIPFlow_1230_io_output_payload_res[65:0];
    _zz_output_payload_res_25 <= multiplierIPFlow_1231_io_output_payload_res[65:0];
    _zz_output_payload_res_26 <= _zz__zz_output_payload_res_26[66:0];
    _zz_output_payload_res_27 <= (_zz__zz_output_payload_res_27 + _zz__zz_output_payload_res_27_3);
    _zz_output_payload_res_28 <= _zz_output_payload_res_19[129:0];
    _zz_output_payload_res_29 <= _zz_output_payload_res_23[129:0];
    _zz_output_payload_res_30 <= _zz__zz_output_payload_res_30[130:0];
    _zz_output_payload_res_31 <= _zz__zz_output_payload_res_31[257:0];
    _zz_io_input_payload_op1_56 <= _zz_io_input_payload_op1_54;
    _zz_io_input_payload_op1_57 <= _zz_io_input_payload_op1_55;
    _zz_io_input_payload_op2_56 <= _zz_io_input_payload_op2_54;
    _zz_io_input_payload_op2_57 <= _zz_io_input_payload_op2_55;
    _zz_io_input_payload_op1_58 <= ({1'b0,_zz_io_input_payload_op1_54} + _zz__zz_io_input_payload_op1_58);
    _zz_io_input_payload_op2_58 <= ({1'b0,_zz_io_input_payload_op2_54} + _zz__zz_io_input_payload_op2_58);
    _zz_io_input_payload_op1_62 <= _zz_io_input_payload_op1_60;
    _zz_io_input_payload_op1_63 <= _zz_io_input_payload_op1_61;
    _zz_io_input_payload_op2_62 <= _zz_io_input_payload_op2_60;
    _zz_io_input_payload_op2_63 <= _zz_io_input_payload_op2_61;
    _zz_io_input_payload_op1_64 <= ({1'b0,_zz_io_input_payload_op1_60} + {1'b0,_zz_io_input_payload_op1_61});
    _zz_io_input_payload_op2_64 <= ({1'b0,_zz_io_input_payload_op2_60} + {1'b0,_zz_io_input_payload_op2_61});
    _zz_output_payload_res_32 <= multiplierIPFlow_1233_io_output_payload_res[65:0];
    _zz_output_payload_res_33 <= multiplierIPFlow_1234_io_output_payload_res[65:0];
    _zz_output_payload_res_34 <= _zz__zz_output_payload_res_34[66:0];
    _zz_output_payload_res_35 <= (_zz__zz_output_payload_res_35 + _zz__zz_output_payload_res_35_3);
    _zz_io_input_payload_op1_68 <= _zz_io_input_payload_op1_66;
    _zz_io_input_payload_op1_69 <= _zz_io_input_payload_op1_67;
    _zz_io_input_payload_op2_68 <= _zz_io_input_payload_op2_66;
    _zz_io_input_payload_op2_69 <= _zz_io_input_payload_op2_67;
    _zz_io_input_payload_op1_70 <= ({1'b0,_zz_io_input_payload_op1_66} + {1'b0,_zz_io_input_payload_op1_67});
    _zz_io_input_payload_op2_70 <= ({1'b0,_zz_io_input_payload_op2_66} + {1'b0,_zz_io_input_payload_op2_67});
    _zz_output_payload_res_36 <= multiplierIPFlow_1236_io_output_payload_res[65:0];
    _zz_output_payload_res_37 <= multiplierIPFlow_1237_io_output_payload_res[65:0];
    _zz_output_payload_res_38 <= _zz__zz_output_payload_res_38[66:0];
    _zz_output_payload_res_39 <= (_zz__zz_output_payload_res_39 + _zz__zz_output_payload_res_39_3);
    _zz_io_input_payload_op1_74 <= _zz_io_input_payload_op1_72;
    _zz_io_input_payload_op1_75 <= _zz_io_input_payload_op1_73;
    _zz_io_input_payload_op2_74 <= _zz_io_input_payload_op2_72;
    _zz_io_input_payload_op2_75 <= _zz_io_input_payload_op2_73;
    _zz_io_input_payload_op1_76 <= ({1'b0,_zz_io_input_payload_op1_72} + {1'b0,_zz_io_input_payload_op1_73});
    _zz_io_input_payload_op2_76 <= ({1'b0,_zz_io_input_payload_op2_72} + {1'b0,_zz_io_input_payload_op2_73});
    _zz_output_payload_res_40 <= multiplierIPFlow_1239_io_output_payload_res[65:0];
    _zz_output_payload_res_41 <= multiplierIPFlow_1240_io_output_payload_res[65:0];
    _zz_output_payload_res_42 <= _zz__zz_output_payload_res_42[66:0];
    _zz_output_payload_res_43 <= (_zz__zz_output_payload_res_43 + _zz__zz_output_payload_res_43_3);
    _zz_output_payload_res_44 <= _zz_output_payload_res_35[129:0];
    _zz_output_payload_res_45 <= _zz_output_payload_res_39[129:0];
    _zz_output_payload_res_46 <= _zz__zz_output_payload_res_46[130:0];
    _zz_output_payload_res_47 <= _zz__zz_output_payload_res_47[257:0];
    _zz_output_payload_res_48 <= _zz_output_payload_res_15[255:0];
    _zz_output_payload_res_49 <= _zz_output_payload_res_31[255:0];
    _zz_output_payload_res_50 <= _zz__zz_output_payload_res_50[256:0];
    output_payload_res <= (_zz_output_payload_res_51 + _zz_output_payload_res_54);
  end


endmodule

module MultiplierFlow (
  input               io_input_valid,
  input      [254:0]  io_input_payload_op1,
  input      [254:0]  io_input_payload_op2,
  output              io_output_valid,
  output     [509:0]  io_output_payload_res,
  input               clk,
  input               resetn
);

  wire       [33:0]   multiplierIPFlow_1215_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1215_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1216_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1216_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1218_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1218_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1219_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1219_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1221_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1221_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1222_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1222_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1224_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1224_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1225_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1225_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1227_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1227_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1228_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1228_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1230_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1230_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1231_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1231_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1233_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1233_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1234_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1234_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1236_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1236_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1237_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1237_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1239_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1239_io_input_payload_op2;
  wire       [33:0]   multiplierIPFlow_1240_io_input_payload_op1;
  wire       [33:0]   multiplierIPFlow_1240_io_input_payload_op2;
  wire                multiplierIPFlow_1215_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1215_io_output_payload_res;
  wire                multiplierIPFlow_1216_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1216_io_output_payload_res;
  wire                multiplierIPFlow_1217_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1217_io_output_payload_res;
  wire                multiplierIPFlow_1218_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1218_io_output_payload_res;
  wire                multiplierIPFlow_1219_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1219_io_output_payload_res;
  wire                multiplierIPFlow_1220_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1220_io_output_payload_res;
  wire                multiplierIPFlow_1221_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1221_io_output_payload_res;
  wire                multiplierIPFlow_1222_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1222_io_output_payload_res;
  wire                multiplierIPFlow_1223_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1223_io_output_payload_res;
  wire                multiplierIPFlow_1224_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1224_io_output_payload_res;
  wire                multiplierIPFlow_1225_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1225_io_output_payload_res;
  wire                multiplierIPFlow_1226_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1226_io_output_payload_res;
  wire                multiplierIPFlow_1227_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1227_io_output_payload_res;
  wire                multiplierIPFlow_1228_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1228_io_output_payload_res;
  wire                multiplierIPFlow_1229_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1229_io_output_payload_res;
  wire                multiplierIPFlow_1230_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1230_io_output_payload_res;
  wire                multiplierIPFlow_1231_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1231_io_output_payload_res;
  wire                multiplierIPFlow_1232_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1232_io_output_payload_res;
  wire                multiplierIPFlow_1233_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1233_io_output_payload_res;
  wire                multiplierIPFlow_1234_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1234_io_output_payload_res;
  wire                multiplierIPFlow_1235_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1235_io_output_payload_res;
  wire                multiplierIPFlow_1236_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1236_io_output_payload_res;
  wire                multiplierIPFlow_1237_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1237_io_output_payload_res;
  wire                multiplierIPFlow_1238_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1238_io_output_payload_res;
  wire                multiplierIPFlow_1239_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1239_io_output_payload_res;
  wire                multiplierIPFlow_1240_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1240_io_output_payload_res;
  wire                multiplierIPFlow_1241_io_output_valid;
  wire       [67:0]   multiplierIPFlow_1241_io_output_payload_res;
  wire       [128:0]  _zz__zz_io_input_payload_op1_4;
  wire       [127:0]  _zz__zz_io_input_payload_op1_4_1;
  wire       [128:0]  _zz__zz_io_input_payload_op2_4;
  wire       [127:0]  _zz__zz_io_input_payload_op2_4_1;
  wire       [65:0]   _zz__zz_io_input_payload_op1_10;
  wire       [64:0]   _zz__zz_io_input_payload_op1_10_1;
  wire       [65:0]   _zz__zz_io_input_payload_op2_10;
  wire       [64:0]   _zz__zz_io_input_payload_op2_10_1;
  wire       [67:0]   _zz__zz_output_payload_res_2;
  wire       [67:0]   _zz__zz_output_payload_res_2_1;
  wire       [131:0]  _zz__zz_output_payload_res_3;
  wire       [131:0]  _zz__zz_output_payload_res_3_1;
  wire       [131:0]  _zz__zz_output_payload_res_3_2;
  wire       [131:0]  _zz__zz_output_payload_res_3_3;
  wire       [99:0]   _zz__zz_output_payload_res_3_4;
  wire       [67:0]   _zz__zz_output_payload_res_6;
  wire       [67:0]   _zz__zz_output_payload_res_6_1;
  wire       [131:0]  _zz__zz_output_payload_res_7;
  wire       [131:0]  _zz__zz_output_payload_res_7_1;
  wire       [131:0]  _zz__zz_output_payload_res_7_2;
  wire       [131:0]  _zz__zz_output_payload_res_7_3;
  wire       [99:0]   _zz__zz_output_payload_res_7_4;
  wire       [67:0]   _zz__zz_output_payload_res_10;
  wire       [67:0]   _zz__zz_output_payload_res_10_1;
  wire       [131:0]  _zz__zz_output_payload_res_11;
  wire       [131:0]  _zz__zz_output_payload_res_11_1;
  wire       [131:0]  _zz__zz_output_payload_res_11_2;
  wire       [131:0]  _zz__zz_output_payload_res_11_3;
  wire       [99:0]   _zz__zz_output_payload_res_11_4;
  wire       [131:0]  _zz__zz_output_payload_res_14;
  wire       [131:0]  _zz__zz_output_payload_res_14_1;
  wire       [259:0]  _zz__zz_output_payload_res_15;
  wire       [259:0]  _zz__zz_output_payload_res_15_1;
  wire       [259:0]  _zz__zz_output_payload_res_15_2;
  wire       [259:0]  _zz__zz_output_payload_res_15_3;
  wire       [259:0]  _zz__zz_output_payload_res_15_4;
  wire       [195:0]  _zz__zz_output_payload_res_15_5;
  wire       [65:0]   _zz__zz_io_input_payload_op1_34;
  wire       [64:0]   _zz__zz_io_input_payload_op1_34_1;
  wire       [65:0]   _zz__zz_io_input_payload_op2_34;
  wire       [64:0]   _zz__zz_io_input_payload_op2_34_1;
  wire       [67:0]   _zz__zz_output_payload_res_18;
  wire       [67:0]   _zz__zz_output_payload_res_18_1;
  wire       [131:0]  _zz__zz_output_payload_res_19;
  wire       [131:0]  _zz__zz_output_payload_res_19_1;
  wire       [131:0]  _zz__zz_output_payload_res_19_2;
  wire       [131:0]  _zz__zz_output_payload_res_19_3;
  wire       [99:0]   _zz__zz_output_payload_res_19_4;
  wire       [67:0]   _zz__zz_output_payload_res_22;
  wire       [67:0]   _zz__zz_output_payload_res_22_1;
  wire       [131:0]  _zz__zz_output_payload_res_23;
  wire       [131:0]  _zz__zz_output_payload_res_23_1;
  wire       [131:0]  _zz__zz_output_payload_res_23_2;
  wire       [131:0]  _zz__zz_output_payload_res_23_3;
  wire       [99:0]   _zz__zz_output_payload_res_23_4;
  wire       [67:0]   _zz__zz_output_payload_res_26;
  wire       [67:0]   _zz__zz_output_payload_res_26_1;
  wire       [131:0]  _zz__zz_output_payload_res_27;
  wire       [131:0]  _zz__zz_output_payload_res_27_1;
  wire       [131:0]  _zz__zz_output_payload_res_27_2;
  wire       [131:0]  _zz__zz_output_payload_res_27_3;
  wire       [99:0]   _zz__zz_output_payload_res_27_4;
  wire       [131:0]  _zz__zz_output_payload_res_30;
  wire       [131:0]  _zz__zz_output_payload_res_30_1;
  wire       [259:0]  _zz__zz_output_payload_res_31;
  wire       [259:0]  _zz__zz_output_payload_res_31_1;
  wire       [259:0]  _zz__zz_output_payload_res_31_2;
  wire       [259:0]  _zz__zz_output_payload_res_31_3;
  wire       [259:0]  _zz__zz_output_payload_res_31_4;
  wire       [195:0]  _zz__zz_output_payload_res_31_5;
  wire       [65:0]   _zz__zz_io_input_payload_op1_58;
  wire       [64:0]   _zz__zz_io_input_payload_op1_58_1;
  wire       [65:0]   _zz__zz_io_input_payload_op2_58;
  wire       [64:0]   _zz__zz_io_input_payload_op2_58_1;
  wire       [67:0]   _zz__zz_output_payload_res_34;
  wire       [67:0]   _zz__zz_output_payload_res_34_1;
  wire       [131:0]  _zz__zz_output_payload_res_35;
  wire       [131:0]  _zz__zz_output_payload_res_35_1;
  wire       [131:0]  _zz__zz_output_payload_res_35_2;
  wire       [131:0]  _zz__zz_output_payload_res_35_3;
  wire       [99:0]   _zz__zz_output_payload_res_35_4;
  wire       [67:0]   _zz__zz_output_payload_res_38;
  wire       [67:0]   _zz__zz_output_payload_res_38_1;
  wire       [131:0]  _zz__zz_output_payload_res_39;
  wire       [131:0]  _zz__zz_output_payload_res_39_1;
  wire       [131:0]  _zz__zz_output_payload_res_39_2;
  wire       [131:0]  _zz__zz_output_payload_res_39_3;
  wire       [99:0]   _zz__zz_output_payload_res_39_4;
  wire       [67:0]   _zz__zz_output_payload_res_42;
  wire       [67:0]   _zz__zz_output_payload_res_42_1;
  wire       [131:0]  _zz__zz_output_payload_res_43;
  wire       [131:0]  _zz__zz_output_payload_res_43_1;
  wire       [131:0]  _zz__zz_output_payload_res_43_2;
  wire       [131:0]  _zz__zz_output_payload_res_43_3;
  wire       [99:0]   _zz__zz_output_payload_res_43_4;
  wire       [131:0]  _zz__zz_output_payload_res_46;
  wire       [131:0]  _zz__zz_output_payload_res_46_1;
  wire       [259:0]  _zz__zz_output_payload_res_47;
  wire       [259:0]  _zz__zz_output_payload_res_47_1;
  wire       [259:0]  _zz__zz_output_payload_res_47_2;
  wire       [259:0]  _zz__zz_output_payload_res_47_3;
  wire       [259:0]  _zz__zz_output_payload_res_47_4;
  wire       [195:0]  _zz__zz_output_payload_res_47_5;
  wire       [257:0]  _zz__zz_output_payload_res_50;
  wire       [257:0]  _zz__zz_output_payload_res_50_1;
  wire       [511:0]  _zz_output_payload_res_51;
  wire       [511:0]  _zz_output_payload_res_52;
  wire       [511:0]  _zz_output_payload_res_53;
  wire       [511:0]  _zz_output_payload_res_54;
  wire       [511:0]  _zz_output_payload_res_55;
  wire       [384:0]  _zz_output_payload_res_56;
  wire       [127:0]  _zz_io_input_payload_op1;
  wire       [126:0]  _zz_io_input_payload_op1_1;
  wire       [127:0]  _zz_io_input_payload_op2;
  wire       [126:0]  _zz_io_input_payload_op2_1;
  reg                 _zz_io_input_valid;
  reg        [127:0]  _zz_io_input_payload_op1_2;
  reg        [126:0]  _zz_io_input_payload_op1_3;
  reg        [127:0]  _zz_io_input_payload_op2_2;
  reg        [126:0]  _zz_io_input_payload_op2_3;
  reg        [128:0]  _zz_io_input_payload_op1_4;
  reg        [128:0]  _zz_io_input_payload_op2_4;
  wire       [128:0]  _zz_io_input_payload_op1_5;
  wire       [128:0]  _zz_io_input_payload_op2_5;
  wire       [64:0]   _zz_io_input_payload_op1_6;
  wire       [63:0]   _zz_io_input_payload_op1_7;
  wire       [64:0]   _zz_io_input_payload_op2_6;
  wire       [63:0]   _zz_io_input_payload_op2_7;
  reg                 _zz_io_input_valid_1;
  reg        [64:0]   _zz_io_input_payload_op1_8;
  reg        [63:0]   _zz_io_input_payload_op1_9;
  reg        [64:0]   _zz_io_input_payload_op2_8;
  reg        [63:0]   _zz_io_input_payload_op2_9;
  reg        [65:0]   _zz_io_input_payload_op1_10;
  reg        [65:0]   _zz_io_input_payload_op2_10;
  wire       [65:0]   _zz_io_input_payload_op1_11;
  wire       [65:0]   _zz_io_input_payload_op2_11;
  wire       [32:0]   _zz_io_input_payload_op1_12;
  wire       [32:0]   _zz_io_input_payload_op1_13;
  wire       [32:0]   _zz_io_input_payload_op2_12;
  wire       [32:0]   _zz_io_input_payload_op2_13;
  reg                 _zz_io_input_valid_2;
  reg        [32:0]   _zz_io_input_payload_op1_14;
  reg        [32:0]   _zz_io_input_payload_op1_15;
  reg        [32:0]   _zz_io_input_payload_op2_14;
  reg        [32:0]   _zz_io_input_payload_op2_15;
  reg        [33:0]   _zz_io_input_payload_op1_16;
  reg        [33:0]   _zz_io_input_payload_op2_16;
  reg                 _zz_output_valid;
  reg        [65:0]   _zz_output_payload_res;
  reg        [65:0]   _zz_output_payload_res_1;
  reg        [66:0]   _zz_output_payload_res_2;
  reg                 _zz_output_valid_1;
  reg        [131:0]  _zz_output_payload_res_3;
  wire       [65:0]   _zz_io_input_payload_op1_17;
  wire       [65:0]   _zz_io_input_payload_op2_17;
  wire       [32:0]   _zz_io_input_payload_op1_18;
  wire       [32:0]   _zz_io_input_payload_op1_19;
  wire       [32:0]   _zz_io_input_payload_op2_18;
  wire       [32:0]   _zz_io_input_payload_op2_19;
  reg                 _zz_io_input_valid_3;
  reg        [32:0]   _zz_io_input_payload_op1_20;
  reg        [32:0]   _zz_io_input_payload_op1_21;
  reg        [32:0]   _zz_io_input_payload_op2_20;
  reg        [32:0]   _zz_io_input_payload_op2_21;
  reg        [33:0]   _zz_io_input_payload_op1_22;
  reg        [33:0]   _zz_io_input_payload_op2_22;
  reg                 _zz_output_valid_2;
  reg        [65:0]   _zz_output_payload_res_4;
  reg        [65:0]   _zz_output_payload_res_5;
  reg        [66:0]   _zz_output_payload_res_6;
  reg                 _zz_output_valid_3;
  reg        [131:0]  _zz_output_payload_res_7;
  wire       [65:0]   _zz_io_input_payload_op1_23;
  wire       [65:0]   _zz_io_input_payload_op2_23;
  wire       [32:0]   _zz_io_input_payload_op1_24;
  wire       [32:0]   _zz_io_input_payload_op1_25;
  wire       [32:0]   _zz_io_input_payload_op2_24;
  wire       [32:0]   _zz_io_input_payload_op2_25;
  reg                 _zz_io_input_valid_4;
  reg        [32:0]   _zz_io_input_payload_op1_26;
  reg        [32:0]   _zz_io_input_payload_op1_27;
  reg        [32:0]   _zz_io_input_payload_op2_26;
  reg        [32:0]   _zz_io_input_payload_op2_27;
  reg        [33:0]   _zz_io_input_payload_op1_28;
  reg        [33:0]   _zz_io_input_payload_op2_28;
  reg                 _zz_output_valid_4;
  reg        [65:0]   _zz_output_payload_res_8;
  reg        [65:0]   _zz_output_payload_res_9;
  reg        [66:0]   _zz_output_payload_res_10;
  reg                 _zz_output_valid_5;
  reg        [131:0]  _zz_output_payload_res_11;
  reg                 _zz_output_valid_6;
  reg        [129:0]  _zz_output_payload_res_12;
  reg        [129:0]  _zz_output_payload_res_13;
  reg        [130:0]  _zz_output_payload_res_14;
  reg                 _zz_output_valid_7;
  reg        [257:0]  _zz_output_payload_res_15;
  wire       [128:0]  _zz_io_input_payload_op1_29;
  wire       [128:0]  _zz_io_input_payload_op2_29;
  wire       [64:0]   _zz_io_input_payload_op1_30;
  wire       [63:0]   _zz_io_input_payload_op1_31;
  wire       [64:0]   _zz_io_input_payload_op2_30;
  wire       [63:0]   _zz_io_input_payload_op2_31;
  reg                 _zz_io_input_valid_5;
  reg        [64:0]   _zz_io_input_payload_op1_32;
  reg        [63:0]   _zz_io_input_payload_op1_33;
  reg        [64:0]   _zz_io_input_payload_op2_32;
  reg        [63:0]   _zz_io_input_payload_op2_33;
  reg        [65:0]   _zz_io_input_payload_op1_34;
  reg        [65:0]   _zz_io_input_payload_op2_34;
  wire       [65:0]   _zz_io_input_payload_op1_35;
  wire       [65:0]   _zz_io_input_payload_op2_35;
  wire       [32:0]   _zz_io_input_payload_op1_36;
  wire       [32:0]   _zz_io_input_payload_op1_37;
  wire       [32:0]   _zz_io_input_payload_op2_36;
  wire       [32:0]   _zz_io_input_payload_op2_37;
  reg                 _zz_io_input_valid_6;
  reg        [32:0]   _zz_io_input_payload_op1_38;
  reg        [32:0]   _zz_io_input_payload_op1_39;
  reg        [32:0]   _zz_io_input_payload_op2_38;
  reg        [32:0]   _zz_io_input_payload_op2_39;
  reg        [33:0]   _zz_io_input_payload_op1_40;
  reg        [33:0]   _zz_io_input_payload_op2_40;
  reg                 _zz_output_valid_8;
  reg        [65:0]   _zz_output_payload_res_16;
  reg        [65:0]   _zz_output_payload_res_17;
  reg        [66:0]   _zz_output_payload_res_18;
  reg                 _zz_output_valid_9;
  reg        [131:0]  _zz_output_payload_res_19;
  wire       [65:0]   _zz_io_input_payload_op1_41;
  wire       [65:0]   _zz_io_input_payload_op2_41;
  wire       [32:0]   _zz_io_input_payload_op1_42;
  wire       [32:0]   _zz_io_input_payload_op1_43;
  wire       [32:0]   _zz_io_input_payload_op2_42;
  wire       [32:0]   _zz_io_input_payload_op2_43;
  reg                 _zz_io_input_valid_7;
  reg        [32:0]   _zz_io_input_payload_op1_44;
  reg        [32:0]   _zz_io_input_payload_op1_45;
  reg        [32:0]   _zz_io_input_payload_op2_44;
  reg        [32:0]   _zz_io_input_payload_op2_45;
  reg        [33:0]   _zz_io_input_payload_op1_46;
  reg        [33:0]   _zz_io_input_payload_op2_46;
  reg                 _zz_output_valid_10;
  reg        [65:0]   _zz_output_payload_res_20;
  reg        [65:0]   _zz_output_payload_res_21;
  reg        [66:0]   _zz_output_payload_res_22;
  reg                 _zz_output_valid_11;
  reg        [131:0]  _zz_output_payload_res_23;
  wire       [65:0]   _zz_io_input_payload_op1_47;
  wire       [65:0]   _zz_io_input_payload_op2_47;
  wire       [32:0]   _zz_io_input_payload_op1_48;
  wire       [32:0]   _zz_io_input_payload_op1_49;
  wire       [32:0]   _zz_io_input_payload_op2_48;
  wire       [32:0]   _zz_io_input_payload_op2_49;
  reg                 _zz_io_input_valid_8;
  reg        [32:0]   _zz_io_input_payload_op1_50;
  reg        [32:0]   _zz_io_input_payload_op1_51;
  reg        [32:0]   _zz_io_input_payload_op2_50;
  reg        [32:0]   _zz_io_input_payload_op2_51;
  reg        [33:0]   _zz_io_input_payload_op1_52;
  reg        [33:0]   _zz_io_input_payload_op2_52;
  reg                 _zz_output_valid_12;
  reg        [65:0]   _zz_output_payload_res_24;
  reg        [65:0]   _zz_output_payload_res_25;
  reg        [66:0]   _zz_output_payload_res_26;
  reg                 _zz_output_valid_13;
  reg        [131:0]  _zz_output_payload_res_27;
  reg                 _zz_output_valid_14;
  reg        [129:0]  _zz_output_payload_res_28;
  reg        [129:0]  _zz_output_payload_res_29;
  reg        [130:0]  _zz_output_payload_res_30;
  reg                 _zz_output_valid_15;
  reg        [257:0]  _zz_output_payload_res_31;
  wire       [128:0]  _zz_io_input_payload_op1_53;
  wire       [128:0]  _zz_io_input_payload_op2_53;
  wire       [64:0]   _zz_io_input_payload_op1_54;
  wire       [63:0]   _zz_io_input_payload_op1_55;
  wire       [64:0]   _zz_io_input_payload_op2_54;
  wire       [63:0]   _zz_io_input_payload_op2_55;
  reg                 _zz_io_input_valid_9;
  reg        [64:0]   _zz_io_input_payload_op1_56;
  reg        [63:0]   _zz_io_input_payload_op1_57;
  reg        [64:0]   _zz_io_input_payload_op2_56;
  reg        [63:0]   _zz_io_input_payload_op2_57;
  reg        [65:0]   _zz_io_input_payload_op1_58;
  reg        [65:0]   _zz_io_input_payload_op2_58;
  wire       [65:0]   _zz_io_input_payload_op1_59;
  wire       [65:0]   _zz_io_input_payload_op2_59;
  wire       [32:0]   _zz_io_input_payload_op1_60;
  wire       [32:0]   _zz_io_input_payload_op1_61;
  wire       [32:0]   _zz_io_input_payload_op2_60;
  wire       [32:0]   _zz_io_input_payload_op2_61;
  reg                 _zz_io_input_valid_10;
  reg        [32:0]   _zz_io_input_payload_op1_62;
  reg        [32:0]   _zz_io_input_payload_op1_63;
  reg        [32:0]   _zz_io_input_payload_op2_62;
  reg        [32:0]   _zz_io_input_payload_op2_63;
  reg        [33:0]   _zz_io_input_payload_op1_64;
  reg        [33:0]   _zz_io_input_payload_op2_64;
  reg                 _zz_output_valid_16;
  reg        [65:0]   _zz_output_payload_res_32;
  reg        [65:0]   _zz_output_payload_res_33;
  reg        [66:0]   _zz_output_payload_res_34;
  reg                 _zz_output_valid_17;
  reg        [131:0]  _zz_output_payload_res_35;
  wire       [65:0]   _zz_io_input_payload_op1_65;
  wire       [65:0]   _zz_io_input_payload_op2_65;
  wire       [32:0]   _zz_io_input_payload_op1_66;
  wire       [32:0]   _zz_io_input_payload_op1_67;
  wire       [32:0]   _zz_io_input_payload_op2_66;
  wire       [32:0]   _zz_io_input_payload_op2_67;
  reg                 _zz_io_input_valid_11;
  reg        [32:0]   _zz_io_input_payload_op1_68;
  reg        [32:0]   _zz_io_input_payload_op1_69;
  reg        [32:0]   _zz_io_input_payload_op2_68;
  reg        [32:0]   _zz_io_input_payload_op2_69;
  reg        [33:0]   _zz_io_input_payload_op1_70;
  reg        [33:0]   _zz_io_input_payload_op2_70;
  reg                 _zz_output_valid_18;
  reg        [65:0]   _zz_output_payload_res_36;
  reg        [65:0]   _zz_output_payload_res_37;
  reg        [66:0]   _zz_output_payload_res_38;
  reg                 _zz_output_valid_19;
  reg        [131:0]  _zz_output_payload_res_39;
  wire       [65:0]   _zz_io_input_payload_op1_71;
  wire       [65:0]   _zz_io_input_payload_op2_71;
  wire       [32:0]   _zz_io_input_payload_op1_72;
  wire       [32:0]   _zz_io_input_payload_op1_73;
  wire       [32:0]   _zz_io_input_payload_op2_72;
  wire       [32:0]   _zz_io_input_payload_op2_73;
  reg                 _zz_io_input_valid_12;
  reg        [32:0]   _zz_io_input_payload_op1_74;
  reg        [32:0]   _zz_io_input_payload_op1_75;
  reg        [32:0]   _zz_io_input_payload_op2_74;
  reg        [32:0]   _zz_io_input_payload_op2_75;
  reg        [33:0]   _zz_io_input_payload_op1_76;
  reg        [33:0]   _zz_io_input_payload_op2_76;
  reg                 _zz_output_valid_20;
  reg        [65:0]   _zz_output_payload_res_40;
  reg        [65:0]   _zz_output_payload_res_41;
  reg        [66:0]   _zz_output_payload_res_42;
  reg                 _zz_output_valid_21;
  reg        [131:0]  _zz_output_payload_res_43;
  reg                 _zz_output_valid_22;
  reg        [129:0]  _zz_output_payload_res_44;
  reg        [129:0]  _zz_output_payload_res_45;
  reg        [130:0]  _zz_output_payload_res_46;
  reg                 _zz_output_valid_23;
  reg        [257:0]  _zz_output_payload_res_47;
  reg                 _zz_output_valid_24;
  reg        [255:0]  _zz_output_payload_res_48;
  reg        [255:0]  _zz_output_payload_res_49;
  reg        [256:0]  _zz_output_payload_res_50;
  reg                 output_valid;
  reg        [509:0]  output_payload_res;

  assign _zz__zz_io_input_payload_op1_4_1 = {1'b0,_zz_io_input_payload_op1_1};
  assign _zz__zz_io_input_payload_op1_4 = {1'd0, _zz__zz_io_input_payload_op1_4_1};
  assign _zz__zz_io_input_payload_op2_4_1 = {1'b0,_zz_io_input_payload_op2_1};
  assign _zz__zz_io_input_payload_op2_4 = {1'd0, _zz__zz_io_input_payload_op2_4_1};
  assign _zz__zz_io_input_payload_op1_10_1 = {1'b0,_zz_io_input_payload_op1_7};
  assign _zz__zz_io_input_payload_op1_10 = {1'd0, _zz__zz_io_input_payload_op1_10_1};
  assign _zz__zz_io_input_payload_op2_10_1 = {1'b0,_zz_io_input_payload_op2_7};
  assign _zz__zz_io_input_payload_op2_10 = {1'd0, _zz__zz_io_input_payload_op2_10_1};
  assign _zz__zz_output_payload_res_2 = (_zz__zz_output_payload_res_2_1 - multiplierIPFlow_1216_io_output_payload_res);
  assign _zz__zz_output_payload_res_2_1 = (multiplierIPFlow_1217_io_output_payload_res - multiplierIPFlow_1215_io_output_payload_res);
  assign _zz__zz_output_payload_res_3 = (_zz__zz_output_payload_res_3_1 + _zz__zz_output_payload_res_3_2);
  assign _zz__zz_output_payload_res_3_1 = ({66'd0,_zz_output_payload_res} <<< 66);
  assign _zz__zz_output_payload_res_3_2 = {66'd0, _zz_output_payload_res_1};
  assign _zz__zz_output_payload_res_3_4 = ({33'd0,_zz_output_payload_res_2} <<< 33);
  assign _zz__zz_output_payload_res_3_3 = {32'd0, _zz__zz_output_payload_res_3_4};
  assign _zz__zz_output_payload_res_6 = (_zz__zz_output_payload_res_6_1 - multiplierIPFlow_1219_io_output_payload_res);
  assign _zz__zz_output_payload_res_6_1 = (multiplierIPFlow_1220_io_output_payload_res - multiplierIPFlow_1218_io_output_payload_res);
  assign _zz__zz_output_payload_res_7 = (_zz__zz_output_payload_res_7_1 + _zz__zz_output_payload_res_7_2);
  assign _zz__zz_output_payload_res_7_1 = ({66'd0,_zz_output_payload_res_4} <<< 66);
  assign _zz__zz_output_payload_res_7_2 = {66'd0, _zz_output_payload_res_5};
  assign _zz__zz_output_payload_res_7_4 = ({33'd0,_zz_output_payload_res_6} <<< 33);
  assign _zz__zz_output_payload_res_7_3 = {32'd0, _zz__zz_output_payload_res_7_4};
  assign _zz__zz_output_payload_res_10 = (_zz__zz_output_payload_res_10_1 - multiplierIPFlow_1222_io_output_payload_res);
  assign _zz__zz_output_payload_res_10_1 = (multiplierIPFlow_1223_io_output_payload_res - multiplierIPFlow_1221_io_output_payload_res);
  assign _zz__zz_output_payload_res_11 = (_zz__zz_output_payload_res_11_1 + _zz__zz_output_payload_res_11_2);
  assign _zz__zz_output_payload_res_11_1 = ({66'd0,_zz_output_payload_res_8} <<< 66);
  assign _zz__zz_output_payload_res_11_2 = {66'd0, _zz_output_payload_res_9};
  assign _zz__zz_output_payload_res_11_4 = ({33'd0,_zz_output_payload_res_10} <<< 33);
  assign _zz__zz_output_payload_res_11_3 = {32'd0, _zz__zz_output_payload_res_11_4};
  assign _zz__zz_output_payload_res_14 = (_zz__zz_output_payload_res_14_1 - _zz_output_payload_res_7);
  assign _zz__zz_output_payload_res_14_1 = (_zz_output_payload_res_11 - _zz_output_payload_res_3);
  assign _zz__zz_output_payload_res_15 = (_zz__zz_output_payload_res_15_1 + _zz__zz_output_payload_res_15_4);
  assign _zz__zz_output_payload_res_15_1 = (_zz__zz_output_payload_res_15_2 + _zz__zz_output_payload_res_15_3);
  assign _zz__zz_output_payload_res_15_2 = ({130'd0,_zz_output_payload_res_12} <<< 130);
  assign _zz__zz_output_payload_res_15_3 = {130'd0, _zz_output_payload_res_13};
  assign _zz__zz_output_payload_res_15_5 = ({65'd0,_zz_output_payload_res_14} <<< 65);
  assign _zz__zz_output_payload_res_15_4 = {64'd0, _zz__zz_output_payload_res_15_5};
  assign _zz__zz_io_input_payload_op1_34_1 = {1'b0,_zz_io_input_payload_op1_31};
  assign _zz__zz_io_input_payload_op1_34 = {1'd0, _zz__zz_io_input_payload_op1_34_1};
  assign _zz__zz_io_input_payload_op2_34_1 = {1'b0,_zz_io_input_payload_op2_31};
  assign _zz__zz_io_input_payload_op2_34 = {1'd0, _zz__zz_io_input_payload_op2_34_1};
  assign _zz__zz_output_payload_res_18 = (_zz__zz_output_payload_res_18_1 - multiplierIPFlow_1225_io_output_payload_res);
  assign _zz__zz_output_payload_res_18_1 = (multiplierIPFlow_1226_io_output_payload_res - multiplierIPFlow_1224_io_output_payload_res);
  assign _zz__zz_output_payload_res_19 = (_zz__zz_output_payload_res_19_1 + _zz__zz_output_payload_res_19_2);
  assign _zz__zz_output_payload_res_19_1 = ({66'd0,_zz_output_payload_res_16} <<< 66);
  assign _zz__zz_output_payload_res_19_2 = {66'd0, _zz_output_payload_res_17};
  assign _zz__zz_output_payload_res_19_4 = ({33'd0,_zz_output_payload_res_18} <<< 33);
  assign _zz__zz_output_payload_res_19_3 = {32'd0, _zz__zz_output_payload_res_19_4};
  assign _zz__zz_output_payload_res_22 = (_zz__zz_output_payload_res_22_1 - multiplierIPFlow_1228_io_output_payload_res);
  assign _zz__zz_output_payload_res_22_1 = (multiplierIPFlow_1229_io_output_payload_res - multiplierIPFlow_1227_io_output_payload_res);
  assign _zz__zz_output_payload_res_23 = (_zz__zz_output_payload_res_23_1 + _zz__zz_output_payload_res_23_2);
  assign _zz__zz_output_payload_res_23_1 = ({66'd0,_zz_output_payload_res_20} <<< 66);
  assign _zz__zz_output_payload_res_23_2 = {66'd0, _zz_output_payload_res_21};
  assign _zz__zz_output_payload_res_23_4 = ({33'd0,_zz_output_payload_res_22} <<< 33);
  assign _zz__zz_output_payload_res_23_3 = {32'd0, _zz__zz_output_payload_res_23_4};
  assign _zz__zz_output_payload_res_26 = (_zz__zz_output_payload_res_26_1 - multiplierIPFlow_1231_io_output_payload_res);
  assign _zz__zz_output_payload_res_26_1 = (multiplierIPFlow_1232_io_output_payload_res - multiplierIPFlow_1230_io_output_payload_res);
  assign _zz__zz_output_payload_res_27 = (_zz__zz_output_payload_res_27_1 + _zz__zz_output_payload_res_27_2);
  assign _zz__zz_output_payload_res_27_1 = ({66'd0,_zz_output_payload_res_24} <<< 66);
  assign _zz__zz_output_payload_res_27_2 = {66'd0, _zz_output_payload_res_25};
  assign _zz__zz_output_payload_res_27_4 = ({33'd0,_zz_output_payload_res_26} <<< 33);
  assign _zz__zz_output_payload_res_27_3 = {32'd0, _zz__zz_output_payload_res_27_4};
  assign _zz__zz_output_payload_res_30 = (_zz__zz_output_payload_res_30_1 - _zz_output_payload_res_23);
  assign _zz__zz_output_payload_res_30_1 = (_zz_output_payload_res_27 - _zz_output_payload_res_19);
  assign _zz__zz_output_payload_res_31 = (_zz__zz_output_payload_res_31_1 + _zz__zz_output_payload_res_31_4);
  assign _zz__zz_output_payload_res_31_1 = (_zz__zz_output_payload_res_31_2 + _zz__zz_output_payload_res_31_3);
  assign _zz__zz_output_payload_res_31_2 = ({130'd0,_zz_output_payload_res_28} <<< 130);
  assign _zz__zz_output_payload_res_31_3 = {130'd0, _zz_output_payload_res_29};
  assign _zz__zz_output_payload_res_31_5 = ({65'd0,_zz_output_payload_res_30} <<< 65);
  assign _zz__zz_output_payload_res_31_4 = {64'd0, _zz__zz_output_payload_res_31_5};
  assign _zz__zz_io_input_payload_op1_58_1 = {1'b0,_zz_io_input_payload_op1_55};
  assign _zz__zz_io_input_payload_op1_58 = {1'd0, _zz__zz_io_input_payload_op1_58_1};
  assign _zz__zz_io_input_payload_op2_58_1 = {1'b0,_zz_io_input_payload_op2_55};
  assign _zz__zz_io_input_payload_op2_58 = {1'd0, _zz__zz_io_input_payload_op2_58_1};
  assign _zz__zz_output_payload_res_34 = (_zz__zz_output_payload_res_34_1 - multiplierIPFlow_1234_io_output_payload_res);
  assign _zz__zz_output_payload_res_34_1 = (multiplierIPFlow_1235_io_output_payload_res - multiplierIPFlow_1233_io_output_payload_res);
  assign _zz__zz_output_payload_res_35 = (_zz__zz_output_payload_res_35_1 + _zz__zz_output_payload_res_35_2);
  assign _zz__zz_output_payload_res_35_1 = ({66'd0,_zz_output_payload_res_32} <<< 66);
  assign _zz__zz_output_payload_res_35_2 = {66'd0, _zz_output_payload_res_33};
  assign _zz__zz_output_payload_res_35_4 = ({33'd0,_zz_output_payload_res_34} <<< 33);
  assign _zz__zz_output_payload_res_35_3 = {32'd0, _zz__zz_output_payload_res_35_4};
  assign _zz__zz_output_payload_res_38 = (_zz__zz_output_payload_res_38_1 - multiplierIPFlow_1237_io_output_payload_res);
  assign _zz__zz_output_payload_res_38_1 = (multiplierIPFlow_1238_io_output_payload_res - multiplierIPFlow_1236_io_output_payload_res);
  assign _zz__zz_output_payload_res_39 = (_zz__zz_output_payload_res_39_1 + _zz__zz_output_payload_res_39_2);
  assign _zz__zz_output_payload_res_39_1 = ({66'd0,_zz_output_payload_res_36} <<< 66);
  assign _zz__zz_output_payload_res_39_2 = {66'd0, _zz_output_payload_res_37};
  assign _zz__zz_output_payload_res_39_4 = ({33'd0,_zz_output_payload_res_38} <<< 33);
  assign _zz__zz_output_payload_res_39_3 = {32'd0, _zz__zz_output_payload_res_39_4};
  assign _zz__zz_output_payload_res_42 = (_zz__zz_output_payload_res_42_1 - multiplierIPFlow_1240_io_output_payload_res);
  assign _zz__zz_output_payload_res_42_1 = (multiplierIPFlow_1241_io_output_payload_res - multiplierIPFlow_1239_io_output_payload_res);
  assign _zz__zz_output_payload_res_43 = (_zz__zz_output_payload_res_43_1 + _zz__zz_output_payload_res_43_2);
  assign _zz__zz_output_payload_res_43_1 = ({66'd0,_zz_output_payload_res_40} <<< 66);
  assign _zz__zz_output_payload_res_43_2 = {66'd0, _zz_output_payload_res_41};
  assign _zz__zz_output_payload_res_43_4 = ({33'd0,_zz_output_payload_res_42} <<< 33);
  assign _zz__zz_output_payload_res_43_3 = {32'd0, _zz__zz_output_payload_res_43_4};
  assign _zz__zz_output_payload_res_46 = (_zz__zz_output_payload_res_46_1 - _zz_output_payload_res_39);
  assign _zz__zz_output_payload_res_46_1 = (_zz_output_payload_res_43 - _zz_output_payload_res_35);
  assign _zz__zz_output_payload_res_47 = (_zz__zz_output_payload_res_47_1 + _zz__zz_output_payload_res_47_4);
  assign _zz__zz_output_payload_res_47_1 = (_zz__zz_output_payload_res_47_2 + _zz__zz_output_payload_res_47_3);
  assign _zz__zz_output_payload_res_47_2 = ({130'd0,_zz_output_payload_res_44} <<< 130);
  assign _zz__zz_output_payload_res_47_3 = {130'd0, _zz_output_payload_res_45};
  assign _zz__zz_output_payload_res_47_5 = ({65'd0,_zz_output_payload_res_46} <<< 65);
  assign _zz__zz_output_payload_res_47_4 = {64'd0, _zz__zz_output_payload_res_47_5};
  assign _zz__zz_output_payload_res_50 = (_zz__zz_output_payload_res_50_1 - _zz_output_payload_res_31);
  assign _zz__zz_output_payload_res_50_1 = (_zz_output_payload_res_47 - _zz_output_payload_res_15);
  assign _zz_output_payload_res_51 = (_zz_output_payload_res_52 + _zz_output_payload_res_55);
  assign _zz_output_payload_res_52 = (_zz_output_payload_res_53 + _zz_output_payload_res_54);
  assign _zz_output_payload_res_53 = ({256'd0,_zz_output_payload_res_48} <<< 256);
  assign _zz_output_payload_res_54 = {256'd0, _zz_output_payload_res_49};
  assign _zz_output_payload_res_56 = ({128'd0,_zz_output_payload_res_50} <<< 128);
  assign _zz_output_payload_res_55 = {127'd0, _zz_output_payload_res_56};
  MultiplierIPFlow multiplierIPFlow_1215 (
    .io_input_valid           (_zz_io_input_valid_2                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1215_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1215_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1215_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1215_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1216 (
    .io_input_valid           (_zz_io_input_valid_2                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1216_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1216_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1216_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1216_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1217 (
    .io_input_valid           (_zz_io_input_valid_2                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_16[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_16[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1217_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1217_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1218 (
    .io_input_valid           (_zz_io_input_valid_3                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1218_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1218_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1218_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1218_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1219 (
    .io_input_valid           (_zz_io_input_valid_3                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1219_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1219_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1219_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1219_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1220 (
    .io_input_valid           (_zz_io_input_valid_3                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_22[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_22[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1220_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1220_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1221 (
    .io_input_valid           (_zz_io_input_valid_4                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1221_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1221_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1221_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1221_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1222 (
    .io_input_valid           (_zz_io_input_valid_4                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1222_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1222_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1222_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1222_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1223 (
    .io_input_valid           (_zz_io_input_valid_4                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_28[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_28[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1223_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1223_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1224 (
    .io_input_valid           (_zz_io_input_valid_6                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1224_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1224_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1224_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1224_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1225 (
    .io_input_valid           (_zz_io_input_valid_6                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1225_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1225_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1225_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1225_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1226 (
    .io_input_valid           (_zz_io_input_valid_6                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_40[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_40[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1226_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1226_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1227 (
    .io_input_valid           (_zz_io_input_valid_7                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1227_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1227_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1227_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1227_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1228 (
    .io_input_valid           (_zz_io_input_valid_7                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1228_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1228_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1228_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1228_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1229 (
    .io_input_valid           (_zz_io_input_valid_7                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_46[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_46[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1229_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1229_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1230 (
    .io_input_valid           (_zz_io_input_valid_8                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1230_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1230_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1230_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1230_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1231 (
    .io_input_valid           (_zz_io_input_valid_8                               ), //i
    .io_input_payload_op1     (multiplierIPFlow_1231_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1231_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1231_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1231_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1232 (
    .io_input_valid           (_zz_io_input_valid_8                               ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_52[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_52[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1232_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1232_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1233 (
    .io_input_valid           (_zz_io_input_valid_10                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1233_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1233_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1233_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1233_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1234 (
    .io_input_valid           (_zz_io_input_valid_10                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1234_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1234_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1234_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1234_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1235 (
    .io_input_valid           (_zz_io_input_valid_10                              ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_64[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_64[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1235_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1235_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1236 (
    .io_input_valid           (_zz_io_input_valid_11                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1236_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1236_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1236_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1236_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1237 (
    .io_input_valid           (_zz_io_input_valid_11                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1237_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1237_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1237_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1237_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1238 (
    .io_input_valid           (_zz_io_input_valid_11                              ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_70[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_70[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1238_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1238_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1239 (
    .io_input_valid           (_zz_io_input_valid_12                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1239_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1239_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1239_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1239_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1240 (
    .io_input_valid           (_zz_io_input_valid_12                              ), //i
    .io_input_payload_op1     (multiplierIPFlow_1240_io_input_payload_op1[33:0]   ), //i
    .io_input_payload_op2     (multiplierIPFlow_1240_io_input_payload_op2[33:0]   ), //i
    .io_output_valid          (multiplierIPFlow_1240_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1240_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  MultiplierIPFlow multiplierIPFlow_1241 (
    .io_input_valid           (_zz_io_input_valid_12                              ), //i
    .io_input_payload_op1     (_zz_io_input_payload_op1_76[33:0]                  ), //i
    .io_input_payload_op2     (_zz_io_input_payload_op2_76[33:0]                  ), //i
    .io_output_valid          (multiplierIPFlow_1241_io_output_valid              ), //o
    .io_output_payload_res    (multiplierIPFlow_1241_io_output_payload_res[67:0]  ), //o
    .clk                      (clk                                                ), //i
    .resetn                   (resetn                                             )  //i
  );
  assign _zz_io_input_payload_op1 = io_input_payload_op1[127 : 0];
  assign _zz_io_input_payload_op1_1 = io_input_payload_op1[254 : 128];
  assign _zz_io_input_payload_op2 = io_input_payload_op2[127 : 0];
  assign _zz_io_input_payload_op2_1 = io_input_payload_op2[254 : 128];
  assign _zz_io_input_payload_op1_5 = {2'd0, _zz_io_input_payload_op1_3};
  assign _zz_io_input_payload_op2_5 = {2'd0, _zz_io_input_payload_op2_3};
  assign _zz_io_input_payload_op1_6 = _zz_io_input_payload_op1_5[64 : 0];
  assign _zz_io_input_payload_op1_7 = _zz_io_input_payload_op1_5[128 : 65];
  assign _zz_io_input_payload_op2_6 = _zz_io_input_payload_op2_5[64 : 0];
  assign _zz_io_input_payload_op2_7 = _zz_io_input_payload_op2_5[128 : 65];
  assign _zz_io_input_payload_op1_11 = {2'd0, _zz_io_input_payload_op1_9};
  assign _zz_io_input_payload_op2_11 = {2'd0, _zz_io_input_payload_op2_9};
  assign _zz_io_input_payload_op1_12 = _zz_io_input_payload_op1_11[32 : 0];
  assign _zz_io_input_payload_op1_13 = _zz_io_input_payload_op1_11[65 : 33];
  assign _zz_io_input_payload_op2_12 = _zz_io_input_payload_op2_11[32 : 0];
  assign _zz_io_input_payload_op2_13 = _zz_io_input_payload_op2_11[65 : 33];
  assign multiplierIPFlow_1215_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_15};
  assign multiplierIPFlow_1215_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_15};
  assign multiplierIPFlow_1216_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_14};
  assign multiplierIPFlow_1216_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_14};
  assign _zz_io_input_payload_op1_17 = {1'd0, _zz_io_input_payload_op1_8};
  assign _zz_io_input_payload_op2_17 = {1'd0, _zz_io_input_payload_op2_8};
  assign _zz_io_input_payload_op1_18 = _zz_io_input_payload_op1_17[32 : 0];
  assign _zz_io_input_payload_op1_19 = _zz_io_input_payload_op1_17[65 : 33];
  assign _zz_io_input_payload_op2_18 = _zz_io_input_payload_op2_17[32 : 0];
  assign _zz_io_input_payload_op2_19 = _zz_io_input_payload_op2_17[65 : 33];
  assign multiplierIPFlow_1218_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_21};
  assign multiplierIPFlow_1218_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_21};
  assign multiplierIPFlow_1219_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_20};
  assign multiplierIPFlow_1219_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_20};
  assign _zz_io_input_payload_op1_23 = _zz_io_input_payload_op1_10;
  assign _zz_io_input_payload_op2_23 = _zz_io_input_payload_op2_10;
  assign _zz_io_input_payload_op1_24 = _zz_io_input_payload_op1_23[32 : 0];
  assign _zz_io_input_payload_op1_25 = _zz_io_input_payload_op1_23[65 : 33];
  assign _zz_io_input_payload_op2_24 = _zz_io_input_payload_op2_23[32 : 0];
  assign _zz_io_input_payload_op2_25 = _zz_io_input_payload_op2_23[65 : 33];
  assign multiplierIPFlow_1221_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_27};
  assign multiplierIPFlow_1221_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_27};
  assign multiplierIPFlow_1222_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_26};
  assign multiplierIPFlow_1222_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_26};
  assign _zz_io_input_payload_op1_29 = {1'd0, _zz_io_input_payload_op1_2};
  assign _zz_io_input_payload_op2_29 = {1'd0, _zz_io_input_payload_op2_2};
  assign _zz_io_input_payload_op1_30 = _zz_io_input_payload_op1_29[64 : 0];
  assign _zz_io_input_payload_op1_31 = _zz_io_input_payload_op1_29[128 : 65];
  assign _zz_io_input_payload_op2_30 = _zz_io_input_payload_op2_29[64 : 0];
  assign _zz_io_input_payload_op2_31 = _zz_io_input_payload_op2_29[128 : 65];
  assign _zz_io_input_payload_op1_35 = {2'd0, _zz_io_input_payload_op1_33};
  assign _zz_io_input_payload_op2_35 = {2'd0, _zz_io_input_payload_op2_33};
  assign _zz_io_input_payload_op1_36 = _zz_io_input_payload_op1_35[32 : 0];
  assign _zz_io_input_payload_op1_37 = _zz_io_input_payload_op1_35[65 : 33];
  assign _zz_io_input_payload_op2_36 = _zz_io_input_payload_op2_35[32 : 0];
  assign _zz_io_input_payload_op2_37 = _zz_io_input_payload_op2_35[65 : 33];
  assign multiplierIPFlow_1224_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_39};
  assign multiplierIPFlow_1224_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_39};
  assign multiplierIPFlow_1225_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_38};
  assign multiplierIPFlow_1225_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_38};
  assign _zz_io_input_payload_op1_41 = {1'd0, _zz_io_input_payload_op1_32};
  assign _zz_io_input_payload_op2_41 = {1'd0, _zz_io_input_payload_op2_32};
  assign _zz_io_input_payload_op1_42 = _zz_io_input_payload_op1_41[32 : 0];
  assign _zz_io_input_payload_op1_43 = _zz_io_input_payload_op1_41[65 : 33];
  assign _zz_io_input_payload_op2_42 = _zz_io_input_payload_op2_41[32 : 0];
  assign _zz_io_input_payload_op2_43 = _zz_io_input_payload_op2_41[65 : 33];
  assign multiplierIPFlow_1227_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_45};
  assign multiplierIPFlow_1227_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_45};
  assign multiplierIPFlow_1228_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_44};
  assign multiplierIPFlow_1228_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_44};
  assign _zz_io_input_payload_op1_47 = _zz_io_input_payload_op1_34;
  assign _zz_io_input_payload_op2_47 = _zz_io_input_payload_op2_34;
  assign _zz_io_input_payload_op1_48 = _zz_io_input_payload_op1_47[32 : 0];
  assign _zz_io_input_payload_op1_49 = _zz_io_input_payload_op1_47[65 : 33];
  assign _zz_io_input_payload_op2_48 = _zz_io_input_payload_op2_47[32 : 0];
  assign _zz_io_input_payload_op2_49 = _zz_io_input_payload_op2_47[65 : 33];
  assign multiplierIPFlow_1230_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_51};
  assign multiplierIPFlow_1230_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_51};
  assign multiplierIPFlow_1231_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_50};
  assign multiplierIPFlow_1231_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_50};
  assign _zz_io_input_payload_op1_53 = _zz_io_input_payload_op1_4;
  assign _zz_io_input_payload_op2_53 = _zz_io_input_payload_op2_4;
  assign _zz_io_input_payload_op1_54 = _zz_io_input_payload_op1_53[64 : 0];
  assign _zz_io_input_payload_op1_55 = _zz_io_input_payload_op1_53[128 : 65];
  assign _zz_io_input_payload_op2_54 = _zz_io_input_payload_op2_53[64 : 0];
  assign _zz_io_input_payload_op2_55 = _zz_io_input_payload_op2_53[128 : 65];
  assign _zz_io_input_payload_op1_59 = {2'd0, _zz_io_input_payload_op1_57};
  assign _zz_io_input_payload_op2_59 = {2'd0, _zz_io_input_payload_op2_57};
  assign _zz_io_input_payload_op1_60 = _zz_io_input_payload_op1_59[32 : 0];
  assign _zz_io_input_payload_op1_61 = _zz_io_input_payload_op1_59[65 : 33];
  assign _zz_io_input_payload_op2_60 = _zz_io_input_payload_op2_59[32 : 0];
  assign _zz_io_input_payload_op2_61 = _zz_io_input_payload_op2_59[65 : 33];
  assign multiplierIPFlow_1233_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_63};
  assign multiplierIPFlow_1233_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_63};
  assign multiplierIPFlow_1234_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_62};
  assign multiplierIPFlow_1234_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_62};
  assign _zz_io_input_payload_op1_65 = {1'd0, _zz_io_input_payload_op1_56};
  assign _zz_io_input_payload_op2_65 = {1'd0, _zz_io_input_payload_op2_56};
  assign _zz_io_input_payload_op1_66 = _zz_io_input_payload_op1_65[32 : 0];
  assign _zz_io_input_payload_op1_67 = _zz_io_input_payload_op1_65[65 : 33];
  assign _zz_io_input_payload_op2_66 = _zz_io_input_payload_op2_65[32 : 0];
  assign _zz_io_input_payload_op2_67 = _zz_io_input_payload_op2_65[65 : 33];
  assign multiplierIPFlow_1236_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_69};
  assign multiplierIPFlow_1236_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_69};
  assign multiplierIPFlow_1237_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_68};
  assign multiplierIPFlow_1237_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_68};
  assign _zz_io_input_payload_op1_71 = _zz_io_input_payload_op1_58;
  assign _zz_io_input_payload_op2_71 = _zz_io_input_payload_op2_58;
  assign _zz_io_input_payload_op1_72 = _zz_io_input_payload_op1_71[32 : 0];
  assign _zz_io_input_payload_op1_73 = _zz_io_input_payload_op1_71[65 : 33];
  assign _zz_io_input_payload_op2_72 = _zz_io_input_payload_op2_71[32 : 0];
  assign _zz_io_input_payload_op2_73 = _zz_io_input_payload_op2_71[65 : 33];
  assign multiplierIPFlow_1239_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_75};
  assign multiplierIPFlow_1239_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_75};
  assign multiplierIPFlow_1240_io_input_payload_op1 = {1'd0, _zz_io_input_payload_op1_74};
  assign multiplierIPFlow_1240_io_input_payload_op2 = {1'd0, _zz_io_input_payload_op2_74};
  assign io_output_valid = output_valid;
  assign io_output_payload_res = output_payload_res;
  always @(posedge clk) begin
    if(!resetn) begin
      _zz_io_input_valid <= 1'b0;
      _zz_io_input_valid_1 <= 1'b0;
      _zz_io_input_valid_2 <= 1'b0;
      _zz_output_valid <= 1'b0;
      _zz_output_valid_1 <= 1'b0;
      _zz_io_input_valid_3 <= 1'b0;
      _zz_output_valid_2 <= 1'b0;
      _zz_output_valid_3 <= 1'b0;
      _zz_io_input_valid_4 <= 1'b0;
      _zz_output_valid_4 <= 1'b0;
      _zz_output_valid_5 <= 1'b0;
      _zz_output_valid_6 <= 1'b0;
      _zz_output_valid_7 <= 1'b0;
      _zz_io_input_valid_5 <= 1'b0;
      _zz_io_input_valid_6 <= 1'b0;
      _zz_output_valid_8 <= 1'b0;
      _zz_output_valid_9 <= 1'b0;
      _zz_io_input_valid_7 <= 1'b0;
      _zz_output_valid_10 <= 1'b0;
      _zz_output_valid_11 <= 1'b0;
      _zz_io_input_valid_8 <= 1'b0;
      _zz_output_valid_12 <= 1'b0;
      _zz_output_valid_13 <= 1'b0;
      _zz_output_valid_14 <= 1'b0;
      _zz_output_valid_15 <= 1'b0;
      _zz_io_input_valid_9 <= 1'b0;
      _zz_io_input_valid_10 <= 1'b0;
      _zz_output_valid_16 <= 1'b0;
      _zz_output_valid_17 <= 1'b0;
      _zz_io_input_valid_11 <= 1'b0;
      _zz_output_valid_18 <= 1'b0;
      _zz_output_valid_19 <= 1'b0;
      _zz_io_input_valid_12 <= 1'b0;
      _zz_output_valid_20 <= 1'b0;
      _zz_output_valid_21 <= 1'b0;
      _zz_output_valid_22 <= 1'b0;
      _zz_output_valid_23 <= 1'b0;
      _zz_output_valid_24 <= 1'b0;
      output_valid <= 1'b0;
    end else begin
      _zz_io_input_valid <= io_input_valid;
      _zz_io_input_valid_1 <= _zz_io_input_valid;
      _zz_io_input_valid_2 <= _zz_io_input_valid_1;
      _zz_output_valid <= ((multiplierIPFlow_1215_io_output_valid && multiplierIPFlow_1216_io_output_valid) && multiplierIPFlow_1217_io_output_valid);
      _zz_output_valid_1 <= _zz_output_valid;
      _zz_io_input_valid_3 <= _zz_io_input_valid_1;
      _zz_output_valid_2 <= ((multiplierIPFlow_1218_io_output_valid && multiplierIPFlow_1219_io_output_valid) && multiplierIPFlow_1220_io_output_valid);
      _zz_output_valid_3 <= _zz_output_valid_2;
      _zz_io_input_valid_4 <= _zz_io_input_valid_1;
      _zz_output_valid_4 <= ((multiplierIPFlow_1221_io_output_valid && multiplierIPFlow_1222_io_output_valid) && multiplierIPFlow_1223_io_output_valid);
      _zz_output_valid_5 <= _zz_output_valid_4;
      _zz_output_valid_6 <= ((_zz_output_valid_1 && _zz_output_valid_3) && _zz_output_valid_5);
      _zz_output_valid_7 <= _zz_output_valid_6;
      _zz_io_input_valid_5 <= _zz_io_input_valid;
      _zz_io_input_valid_6 <= _zz_io_input_valid_5;
      _zz_output_valid_8 <= ((multiplierIPFlow_1224_io_output_valid && multiplierIPFlow_1225_io_output_valid) && multiplierIPFlow_1226_io_output_valid);
      _zz_output_valid_9 <= _zz_output_valid_8;
      _zz_io_input_valid_7 <= _zz_io_input_valid_5;
      _zz_output_valid_10 <= ((multiplierIPFlow_1227_io_output_valid && multiplierIPFlow_1228_io_output_valid) && multiplierIPFlow_1229_io_output_valid);
      _zz_output_valid_11 <= _zz_output_valid_10;
      _zz_io_input_valid_8 <= _zz_io_input_valid_5;
      _zz_output_valid_12 <= ((multiplierIPFlow_1230_io_output_valid && multiplierIPFlow_1231_io_output_valid) && multiplierIPFlow_1232_io_output_valid);
      _zz_output_valid_13 <= _zz_output_valid_12;
      _zz_output_valid_14 <= ((_zz_output_valid_9 && _zz_output_valid_11) && _zz_output_valid_13);
      _zz_output_valid_15 <= _zz_output_valid_14;
      _zz_io_input_valid_9 <= _zz_io_input_valid;
      _zz_io_input_valid_10 <= _zz_io_input_valid_9;
      _zz_output_valid_16 <= ((multiplierIPFlow_1233_io_output_valid && multiplierIPFlow_1234_io_output_valid) && multiplierIPFlow_1235_io_output_valid);
      _zz_output_valid_17 <= _zz_output_valid_16;
      _zz_io_input_valid_11 <= _zz_io_input_valid_9;
      _zz_output_valid_18 <= ((multiplierIPFlow_1236_io_output_valid && multiplierIPFlow_1237_io_output_valid) && multiplierIPFlow_1238_io_output_valid);
      _zz_output_valid_19 <= _zz_output_valid_18;
      _zz_io_input_valid_12 <= _zz_io_input_valid_9;
      _zz_output_valid_20 <= ((multiplierIPFlow_1239_io_output_valid && multiplierIPFlow_1240_io_output_valid) && multiplierIPFlow_1241_io_output_valid);
      _zz_output_valid_21 <= _zz_output_valid_20;
      _zz_output_valid_22 <= ((_zz_output_valid_17 && _zz_output_valid_19) && _zz_output_valid_21);
      _zz_output_valid_23 <= _zz_output_valid_22;
      _zz_output_valid_24 <= ((_zz_output_valid_7 && _zz_output_valid_15) && _zz_output_valid_23);
      output_valid <= _zz_output_valid_24;
    end
  end

  always @(posedge clk) begin
    _zz_io_input_payload_op1_2 <= _zz_io_input_payload_op1;
    _zz_io_input_payload_op1_3 <= _zz_io_input_payload_op1_1;
    _zz_io_input_payload_op2_2 <= _zz_io_input_payload_op2;
    _zz_io_input_payload_op2_3 <= _zz_io_input_payload_op2_1;
    _zz_io_input_payload_op1_4 <= ({1'b0,_zz_io_input_payload_op1} + _zz__zz_io_input_payload_op1_4);
    _zz_io_input_payload_op2_4 <= ({1'b0,_zz_io_input_payload_op2} + _zz__zz_io_input_payload_op2_4);
    _zz_io_input_payload_op1_8 <= _zz_io_input_payload_op1_6;
    _zz_io_input_payload_op1_9 <= _zz_io_input_payload_op1_7;
    _zz_io_input_payload_op2_8 <= _zz_io_input_payload_op2_6;
    _zz_io_input_payload_op2_9 <= _zz_io_input_payload_op2_7;
    _zz_io_input_payload_op1_10 <= ({1'b0,_zz_io_input_payload_op1_6} + _zz__zz_io_input_payload_op1_10);
    _zz_io_input_payload_op2_10 <= ({1'b0,_zz_io_input_payload_op2_6} + _zz__zz_io_input_payload_op2_10);
    _zz_io_input_payload_op1_14 <= _zz_io_input_payload_op1_12;
    _zz_io_input_payload_op1_15 <= _zz_io_input_payload_op1_13;
    _zz_io_input_payload_op2_14 <= _zz_io_input_payload_op2_12;
    _zz_io_input_payload_op2_15 <= _zz_io_input_payload_op2_13;
    _zz_io_input_payload_op1_16 <= ({1'b0,_zz_io_input_payload_op1_12} + {1'b0,_zz_io_input_payload_op1_13});
    _zz_io_input_payload_op2_16 <= ({1'b0,_zz_io_input_payload_op2_12} + {1'b0,_zz_io_input_payload_op2_13});
    _zz_output_payload_res <= multiplierIPFlow_1215_io_output_payload_res[65:0];
    _zz_output_payload_res_1 <= multiplierIPFlow_1216_io_output_payload_res[65:0];
    _zz_output_payload_res_2 <= _zz__zz_output_payload_res_2[66:0];
    _zz_output_payload_res_3 <= (_zz__zz_output_payload_res_3 + _zz__zz_output_payload_res_3_3);
    _zz_io_input_payload_op1_20 <= _zz_io_input_payload_op1_18;
    _zz_io_input_payload_op1_21 <= _zz_io_input_payload_op1_19;
    _zz_io_input_payload_op2_20 <= _zz_io_input_payload_op2_18;
    _zz_io_input_payload_op2_21 <= _zz_io_input_payload_op2_19;
    _zz_io_input_payload_op1_22 <= ({1'b0,_zz_io_input_payload_op1_18} + {1'b0,_zz_io_input_payload_op1_19});
    _zz_io_input_payload_op2_22 <= ({1'b0,_zz_io_input_payload_op2_18} + {1'b0,_zz_io_input_payload_op2_19});
    _zz_output_payload_res_4 <= multiplierIPFlow_1218_io_output_payload_res[65:0];
    _zz_output_payload_res_5 <= multiplierIPFlow_1219_io_output_payload_res[65:0];
    _zz_output_payload_res_6 <= _zz__zz_output_payload_res_6[66:0];
    _zz_output_payload_res_7 <= (_zz__zz_output_payload_res_7 + _zz__zz_output_payload_res_7_3);
    _zz_io_input_payload_op1_26 <= _zz_io_input_payload_op1_24;
    _zz_io_input_payload_op1_27 <= _zz_io_input_payload_op1_25;
    _zz_io_input_payload_op2_26 <= _zz_io_input_payload_op2_24;
    _zz_io_input_payload_op2_27 <= _zz_io_input_payload_op2_25;
    _zz_io_input_payload_op1_28 <= ({1'b0,_zz_io_input_payload_op1_24} + {1'b0,_zz_io_input_payload_op1_25});
    _zz_io_input_payload_op2_28 <= ({1'b0,_zz_io_input_payload_op2_24} + {1'b0,_zz_io_input_payload_op2_25});
    _zz_output_payload_res_8 <= multiplierIPFlow_1221_io_output_payload_res[65:0];
    _zz_output_payload_res_9 <= multiplierIPFlow_1222_io_output_payload_res[65:0];
    _zz_output_payload_res_10 <= _zz__zz_output_payload_res_10[66:0];
    _zz_output_payload_res_11 <= (_zz__zz_output_payload_res_11 + _zz__zz_output_payload_res_11_3);
    _zz_output_payload_res_12 <= _zz_output_payload_res_3[129:0];
    _zz_output_payload_res_13 <= _zz_output_payload_res_7[129:0];
    _zz_output_payload_res_14 <= _zz__zz_output_payload_res_14[130:0];
    _zz_output_payload_res_15 <= _zz__zz_output_payload_res_15[257:0];
    _zz_io_input_payload_op1_32 <= _zz_io_input_payload_op1_30;
    _zz_io_input_payload_op1_33 <= _zz_io_input_payload_op1_31;
    _zz_io_input_payload_op2_32 <= _zz_io_input_payload_op2_30;
    _zz_io_input_payload_op2_33 <= _zz_io_input_payload_op2_31;
    _zz_io_input_payload_op1_34 <= ({1'b0,_zz_io_input_payload_op1_30} + _zz__zz_io_input_payload_op1_34);
    _zz_io_input_payload_op2_34 <= ({1'b0,_zz_io_input_payload_op2_30} + _zz__zz_io_input_payload_op2_34);
    _zz_io_input_payload_op1_38 <= _zz_io_input_payload_op1_36;
    _zz_io_input_payload_op1_39 <= _zz_io_input_payload_op1_37;
    _zz_io_input_payload_op2_38 <= _zz_io_input_payload_op2_36;
    _zz_io_input_payload_op2_39 <= _zz_io_input_payload_op2_37;
    _zz_io_input_payload_op1_40 <= ({1'b0,_zz_io_input_payload_op1_36} + {1'b0,_zz_io_input_payload_op1_37});
    _zz_io_input_payload_op2_40 <= ({1'b0,_zz_io_input_payload_op2_36} + {1'b0,_zz_io_input_payload_op2_37});
    _zz_output_payload_res_16 <= multiplierIPFlow_1224_io_output_payload_res[65:0];
    _zz_output_payload_res_17 <= multiplierIPFlow_1225_io_output_payload_res[65:0];
    _zz_output_payload_res_18 <= _zz__zz_output_payload_res_18[66:0];
    _zz_output_payload_res_19 <= (_zz__zz_output_payload_res_19 + _zz__zz_output_payload_res_19_3);
    _zz_io_input_payload_op1_44 <= _zz_io_input_payload_op1_42;
    _zz_io_input_payload_op1_45 <= _zz_io_input_payload_op1_43;
    _zz_io_input_payload_op2_44 <= _zz_io_input_payload_op2_42;
    _zz_io_input_payload_op2_45 <= _zz_io_input_payload_op2_43;
    _zz_io_input_payload_op1_46 <= ({1'b0,_zz_io_input_payload_op1_42} + {1'b0,_zz_io_input_payload_op1_43});
    _zz_io_input_payload_op2_46 <= ({1'b0,_zz_io_input_payload_op2_42} + {1'b0,_zz_io_input_payload_op2_43});
    _zz_output_payload_res_20 <= multiplierIPFlow_1227_io_output_payload_res[65:0];
    _zz_output_payload_res_21 <= multiplierIPFlow_1228_io_output_payload_res[65:0];
    _zz_output_payload_res_22 <= _zz__zz_output_payload_res_22[66:0];
    _zz_output_payload_res_23 <= (_zz__zz_output_payload_res_23 + _zz__zz_output_payload_res_23_3);
    _zz_io_input_payload_op1_50 <= _zz_io_input_payload_op1_48;
    _zz_io_input_payload_op1_51 <= _zz_io_input_payload_op1_49;
    _zz_io_input_payload_op2_50 <= _zz_io_input_payload_op2_48;
    _zz_io_input_payload_op2_51 <= _zz_io_input_payload_op2_49;
    _zz_io_input_payload_op1_52 <= ({1'b0,_zz_io_input_payload_op1_48} + {1'b0,_zz_io_input_payload_op1_49});
    _zz_io_input_payload_op2_52 <= ({1'b0,_zz_io_input_payload_op2_48} + {1'b0,_zz_io_input_payload_op2_49});
    _zz_output_payload_res_24 <= multiplierIPFlow_1230_io_output_payload_res[65:0];
    _zz_output_payload_res_25 <= multiplierIPFlow_1231_io_output_payload_res[65:0];
    _zz_output_payload_res_26 <= _zz__zz_output_payload_res_26[66:0];
    _zz_output_payload_res_27 <= (_zz__zz_output_payload_res_27 + _zz__zz_output_payload_res_27_3);
    _zz_output_payload_res_28 <= _zz_output_payload_res_19[129:0];
    _zz_output_payload_res_29 <= _zz_output_payload_res_23[129:0];
    _zz_output_payload_res_30 <= _zz__zz_output_payload_res_30[130:0];
    _zz_output_payload_res_31 <= _zz__zz_output_payload_res_31[257:0];
    _zz_io_input_payload_op1_56 <= _zz_io_input_payload_op1_54;
    _zz_io_input_payload_op1_57 <= _zz_io_input_payload_op1_55;
    _zz_io_input_payload_op2_56 <= _zz_io_input_payload_op2_54;
    _zz_io_input_payload_op2_57 <= _zz_io_input_payload_op2_55;
    _zz_io_input_payload_op1_58 <= ({1'b0,_zz_io_input_payload_op1_54} + _zz__zz_io_input_payload_op1_58);
    _zz_io_input_payload_op2_58 <= ({1'b0,_zz_io_input_payload_op2_54} + _zz__zz_io_input_payload_op2_58);
    _zz_io_input_payload_op1_62 <= _zz_io_input_payload_op1_60;
    _zz_io_input_payload_op1_63 <= _zz_io_input_payload_op1_61;
    _zz_io_input_payload_op2_62 <= _zz_io_input_payload_op2_60;
    _zz_io_input_payload_op2_63 <= _zz_io_input_payload_op2_61;
    _zz_io_input_payload_op1_64 <= ({1'b0,_zz_io_input_payload_op1_60} + {1'b0,_zz_io_input_payload_op1_61});
    _zz_io_input_payload_op2_64 <= ({1'b0,_zz_io_input_payload_op2_60} + {1'b0,_zz_io_input_payload_op2_61});
    _zz_output_payload_res_32 <= multiplierIPFlow_1233_io_output_payload_res[65:0];
    _zz_output_payload_res_33 <= multiplierIPFlow_1234_io_output_payload_res[65:0];
    _zz_output_payload_res_34 <= _zz__zz_output_payload_res_34[66:0];
    _zz_output_payload_res_35 <= (_zz__zz_output_payload_res_35 + _zz__zz_output_payload_res_35_3);
    _zz_io_input_payload_op1_68 <= _zz_io_input_payload_op1_66;
    _zz_io_input_payload_op1_69 <= _zz_io_input_payload_op1_67;
    _zz_io_input_payload_op2_68 <= _zz_io_input_payload_op2_66;
    _zz_io_input_payload_op2_69 <= _zz_io_input_payload_op2_67;
    _zz_io_input_payload_op1_70 <= ({1'b0,_zz_io_input_payload_op1_66} + {1'b0,_zz_io_input_payload_op1_67});
    _zz_io_input_payload_op2_70 <= ({1'b0,_zz_io_input_payload_op2_66} + {1'b0,_zz_io_input_payload_op2_67});
    _zz_output_payload_res_36 <= multiplierIPFlow_1236_io_output_payload_res[65:0];
    _zz_output_payload_res_37 <= multiplierIPFlow_1237_io_output_payload_res[65:0];
    _zz_output_payload_res_38 <= _zz__zz_output_payload_res_38[66:0];
    _zz_output_payload_res_39 <= (_zz__zz_output_payload_res_39 + _zz__zz_output_payload_res_39_3);
    _zz_io_input_payload_op1_74 <= _zz_io_input_payload_op1_72;
    _zz_io_input_payload_op1_75 <= _zz_io_input_payload_op1_73;
    _zz_io_input_payload_op2_74 <= _zz_io_input_payload_op2_72;
    _zz_io_input_payload_op2_75 <= _zz_io_input_payload_op2_73;
    _zz_io_input_payload_op1_76 <= ({1'b0,_zz_io_input_payload_op1_72} + {1'b0,_zz_io_input_payload_op1_73});
    _zz_io_input_payload_op2_76 <= ({1'b0,_zz_io_input_payload_op2_72} + {1'b0,_zz_io_input_payload_op2_73});
    _zz_output_payload_res_40 <= multiplierIPFlow_1239_io_output_payload_res[65:0];
    _zz_output_payload_res_41 <= multiplierIPFlow_1240_io_output_payload_res[65:0];
    _zz_output_payload_res_42 <= _zz__zz_output_payload_res_42[66:0];
    _zz_output_payload_res_43 <= (_zz__zz_output_payload_res_43 + _zz__zz_output_payload_res_43_3);
    _zz_output_payload_res_44 <= _zz_output_payload_res_35[129:0];
    _zz_output_payload_res_45 <= _zz_output_payload_res_39[129:0];
    _zz_output_payload_res_46 <= _zz__zz_output_payload_res_46[130:0];
    _zz_output_payload_res_47 <= _zz__zz_output_payload_res_47[257:0];
    _zz_output_payload_res_48 <= _zz_output_payload_res_15[255:0];
    _zz_output_payload_res_49 <= _zz_output_payload_res_31[255:0];
    _zz_output_payload_res_50 <= _zz__zz_output_payload_res_50[256:0];
    output_payload_res <= _zz_output_payload_res_51[509:0];
  end


endmodule

module MatrixConstantMem_13 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  output     [254:0]  io_data_9,
  output     [254:0]  io_data_10,
  output     [254:0]  io_data_11,
  input      [5:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  reg        [254:0]  _zz_mdsMem_5_port0;
  reg        [254:0]  _zz_mdsMem_6_port0;
  reg        [254:0]  _zz_mdsMem_7_port0;
  reg        [254:0]  _zz_mdsMem_8_port0;
  reg        [254:0]  _zz_mdsMem_9_port0;
  reg        [254:0]  _zz_mdsMem_10_port0;
  reg        [254:0]  _zz_mdsMem_11_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire                _zz_mdsMem_5_port;
  wire                _zz_io_data_5;
  wire                _zz_mdsMem_6_port;
  wire                _zz_io_data_6;
  wire                _zz_mdsMem_7_port;
  wire                _zz_io_data_7;
  wire                _zz_mdsMem_8_port;
  wire                _zz_io_data_8;
  wire                _zz_mdsMem_9_port;
  wire                _zz_io_data_9;
  wire                _zz_mdsMem_10_port;
  wire                _zz_io_data_10;
  wire                _zz_mdsMem_11_port;
  wire                _zz_io_data_11;
  wire       [254:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [254:0]  mdsMatrix_0_2;
  wire       [253:0]  mdsMatrix_0_3;
  wire       [253:0]  mdsMatrix_0_4;
  wire       [253:0]  mdsMatrix_0_5;
  wire       [251:0]  mdsMatrix_0_6;
  wire       [254:0]  mdsMatrix_0_7;
  wire       [254:0]  mdsMatrix_0_8;
  wire       [252:0]  mdsMatrix_0_9;
  wire       [253:0]  mdsMatrix_0_10;
  wire       [253:0]  mdsMatrix_0_11;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [253:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [254:0]  mdsMatrix_1_3;
  wire       [250:0]  mdsMatrix_1_4;
  wire       [254:0]  mdsMatrix_1_5;
  wire       [254:0]  mdsMatrix_1_6;
  wire       [252:0]  mdsMatrix_1_7;
  wire       [254:0]  mdsMatrix_1_8;
  wire       [254:0]  mdsMatrix_1_9;
  wire       [249:0]  mdsMatrix_1_10;
  wire       [252:0]  mdsMatrix_1_11;
  wire       [254:0]  mdsMatrix_2_0;
  wire       [252:0]  mdsMatrix_2_1;
  wire       [253:0]  mdsMatrix_2_2;
  wire       [253:0]  mdsMatrix_2_3;
  wire       [253:0]  mdsMatrix_2_4;
  wire       [252:0]  mdsMatrix_2_5;
  wire       [254:0]  mdsMatrix_2_6;
  wire       [252:0]  mdsMatrix_2_7;
  wire       [251:0]  mdsMatrix_2_8;
  wire       [249:0]  mdsMatrix_2_9;
  wire       [251:0]  mdsMatrix_2_10;
  wire       [254:0]  mdsMatrix_2_11;
  wire       [254:0]  mdsMatrix_3_0;
  wire       [252:0]  mdsMatrix_3_1;
  wire       [253:0]  mdsMatrix_3_2;
  wire       [254:0]  mdsMatrix_3_3;
  wire       [254:0]  mdsMatrix_3_4;
  wire       [253:0]  mdsMatrix_3_5;
  wire       [253:0]  mdsMatrix_3_6;
  wire       [251:0]  mdsMatrix_3_7;
  wire       [253:0]  mdsMatrix_3_8;
  wire       [254:0]  mdsMatrix_3_9;
  wire       [254:0]  mdsMatrix_3_10;
  wire       [254:0]  mdsMatrix_3_11;
  wire       [254:0]  mdsMatrix_4_0;
  wire       [252:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [252:0]  mdsMatrix_4_3;
  wire       [253:0]  mdsMatrix_4_4;
  wire       [251:0]  mdsMatrix_4_5;
  wire       [252:0]  mdsMatrix_4_6;
  wire       [254:0]  mdsMatrix_4_7;
  wire       [254:0]  mdsMatrix_4_8;
  wire       [252:0]  mdsMatrix_4_9;
  wire       [251:0]  mdsMatrix_4_10;
  wire       [254:0]  mdsMatrix_4_11;
  wire       [254:0]  mdsMatrix_5_0;
  wire       [254:0]  mdsMatrix_5_1;
  wire       [254:0]  mdsMatrix_5_2;
  wire       [253:0]  mdsMatrix_5_3;
  wire       [252:0]  mdsMatrix_5_4;
  wire       [254:0]  mdsMatrix_5_5;
  wire       [251:0]  mdsMatrix_5_6;
  wire       [249:0]  mdsMatrix_5_7;
  wire       [247:0]  mdsMatrix_5_8;
  wire       [253:0]  mdsMatrix_5_9;
  wire       [254:0]  mdsMatrix_5_10;
  wire       [253:0]  mdsMatrix_5_11;
  wire       [254:0]  mdsMatrix_6_0;
  wire       [254:0]  mdsMatrix_6_1;
  wire       [251:0]  mdsMatrix_6_2;
  wire       [253:0]  mdsMatrix_6_3;
  wire       [254:0]  mdsMatrix_6_4;
  wire       [252:0]  mdsMatrix_6_5;
  wire       [253:0]  mdsMatrix_6_6;
  wire       [249:0]  mdsMatrix_6_7;
  wire       [254:0]  mdsMatrix_6_8;
  wire       [251:0]  mdsMatrix_6_9;
  wire       [250:0]  mdsMatrix_6_10;
  wire       [253:0]  mdsMatrix_6_11;
  wire       [254:0]  mdsMatrix_7_0;
  wire       [252:0]  mdsMatrix_7_1;
  wire       [253:0]  mdsMatrix_7_2;
  wire       [253:0]  mdsMatrix_7_3;
  wire       [254:0]  mdsMatrix_7_4;
  wire       [253:0]  mdsMatrix_7_5;
  wire       [253:0]  mdsMatrix_7_6;
  wire       [254:0]  mdsMatrix_7_7;
  wire       [254:0]  mdsMatrix_7_8;
  wire       [253:0]  mdsMatrix_7_9;
  wire       [253:0]  mdsMatrix_7_10;
  wire       [253:0]  mdsMatrix_7_11;
  wire       [254:0]  mdsMatrix_8_0;
  wire       [254:0]  mdsMatrix_8_1;
  wire       [254:0]  mdsMatrix_8_2;
  wire       [254:0]  mdsMatrix_8_3;
  wire       [253:0]  mdsMatrix_8_4;
  wire       [254:0]  mdsMatrix_8_5;
  wire       [254:0]  mdsMatrix_8_6;
  wire       [248:0]  mdsMatrix_8_7;
  wire       [252:0]  mdsMatrix_8_8;
  wire       [251:0]  mdsMatrix_8_9;
  wire       [253:0]  mdsMatrix_8_10;
  wire       [253:0]  mdsMatrix_8_11;
  wire       [254:0]  mdsMatrix_9_0;
  wire       [252:0]  mdsMatrix_9_1;
  wire       [253:0]  mdsMatrix_9_2;
  wire       [254:0]  mdsMatrix_9_3;
  wire       [253:0]  mdsMatrix_9_4;
  wire       [252:0]  mdsMatrix_9_5;
  wire       [254:0]  mdsMatrix_9_6;
  wire       [253:0]  mdsMatrix_9_7;
  wire       [252:0]  mdsMatrix_9_8;
  wire       [252:0]  mdsMatrix_9_9;
  wire       [253:0]  mdsMatrix_9_10;
  wire       [254:0]  mdsMatrix_9_11;
  wire       [254:0]  mdsMatrix_10_0;
  wire       [254:0]  mdsMatrix_10_1;
  wire       [254:0]  mdsMatrix_10_2;
  wire       [254:0]  mdsMatrix_10_3;
  wire       [251:0]  mdsMatrix_10_4;
  wire       [254:0]  mdsMatrix_10_5;
  wire       [252:0]  mdsMatrix_10_6;
  wire       [253:0]  mdsMatrix_10_7;
  wire       [254:0]  mdsMatrix_10_8;
  wire       [253:0]  mdsMatrix_10_9;
  wire       [252:0]  mdsMatrix_10_10;
  wire       [254:0]  mdsMatrix_10_11;
  wire       [254:0]  mdsMatrix_11_0;
  wire       [253:0]  mdsMatrix_11_1;
  wire       [251:0]  mdsMatrix_11_2;
  wire       [254:0]  mdsMatrix_11_3;
  wire       [254:0]  mdsMatrix_11_4;
  wire       [254:0]  mdsMatrix_11_5;
  wire       [252:0]  mdsMatrix_11_6;
  wire       [254:0]  mdsMatrix_11_7;
  wire       [252:0]  mdsMatrix_11_8;
  wire       [252:0]  mdsMatrix_11_9;
  wire       [253:0]  mdsMatrix_11_10;
  wire       [253:0]  mdsMatrix_11_11;
  wire       [254:0]  mdsMatrix_12_0;
  wire       [254:0]  mdsMatrix_12_1;
  wire       [254:0]  mdsMatrix_12_2;
  wire       [254:0]  mdsMatrix_12_3;
  wire       [252:0]  mdsMatrix_12_4;
  wire       [253:0]  mdsMatrix_12_5;
  wire       [254:0]  mdsMatrix_12_6;
  wire       [253:0]  mdsMatrix_12_7;
  wire       [254:0]  mdsMatrix_12_8;
  wire       [252:0]  mdsMatrix_12_9;
  wire       [254:0]  mdsMatrix_12_10;
  wire       [254:0]  mdsMatrix_12_11;
  wire       [254:0]  mdsMatrix_13_0;
  wire       [254:0]  mdsMatrix_13_1;
  wire       [254:0]  mdsMatrix_13_2;
  wire       [254:0]  mdsMatrix_13_3;
  wire       [251:0]  mdsMatrix_13_4;
  wire       [254:0]  mdsMatrix_13_5;
  wire       [252:0]  mdsMatrix_13_6;
  wire       [249:0]  mdsMatrix_13_7;
  wire       [252:0]  mdsMatrix_13_8;
  wire       [254:0]  mdsMatrix_13_9;
  wire       [254:0]  mdsMatrix_13_10;
  wire       [253:0]  mdsMatrix_13_11;
  wire       [254:0]  mdsMatrix_14_0;
  wire       [254:0]  mdsMatrix_14_1;
  wire       [252:0]  mdsMatrix_14_2;
  wire       [253:0]  mdsMatrix_14_3;
  wire       [251:0]  mdsMatrix_14_4;
  wire       [252:0]  mdsMatrix_14_5;
  wire       [254:0]  mdsMatrix_14_6;
  wire       [254:0]  mdsMatrix_14_7;
  wire       [254:0]  mdsMatrix_14_8;
  wire       [254:0]  mdsMatrix_14_9;
  wire       [254:0]  mdsMatrix_14_10;
  wire       [253:0]  mdsMatrix_14_11;
  wire       [254:0]  mdsMatrix_15_0;
  wire       [252:0]  mdsMatrix_15_1;
  wire       [253:0]  mdsMatrix_15_2;
  wire       [253:0]  mdsMatrix_15_3;
  wire       [252:0]  mdsMatrix_15_4;
  wire       [254:0]  mdsMatrix_15_5;
  wire       [254:0]  mdsMatrix_15_6;
  wire       [252:0]  mdsMatrix_15_7;
  wire       [252:0]  mdsMatrix_15_8;
  wire       [254:0]  mdsMatrix_15_9;
  wire       [254:0]  mdsMatrix_15_10;
  wire       [254:0]  mdsMatrix_15_11;
  wire       [254:0]  mdsMatrix_16_0;
  wire       [254:0]  mdsMatrix_16_1;
  wire       [253:0]  mdsMatrix_16_2;
  wire       [254:0]  mdsMatrix_16_3;
  wire       [251:0]  mdsMatrix_16_4;
  wire       [253:0]  mdsMatrix_16_5;
  wire       [253:0]  mdsMatrix_16_6;
  wire       [252:0]  mdsMatrix_16_7;
  wire       [252:0]  mdsMatrix_16_8;
  wire       [246:0]  mdsMatrix_16_9;
  wire       [254:0]  mdsMatrix_16_10;
  wire       [253:0]  mdsMatrix_16_11;
  wire       [254:0]  mdsMatrix_17_0;
  wire       [250:0]  mdsMatrix_17_1;
  wire       [254:0]  mdsMatrix_17_2;
  wire       [253:0]  mdsMatrix_17_3;
  wire       [252:0]  mdsMatrix_17_4;
  wire       [253:0]  mdsMatrix_17_5;
  wire       [254:0]  mdsMatrix_17_6;
  wire       [254:0]  mdsMatrix_17_7;
  wire       [254:0]  mdsMatrix_17_8;
  wire       [254:0]  mdsMatrix_17_9;
  wire       [253:0]  mdsMatrix_17_10;
  wire       [251:0]  mdsMatrix_17_11;
  wire       [254:0]  mdsMatrix_18_0;
  wire       [252:0]  mdsMatrix_18_1;
  wire       [251:0]  mdsMatrix_18_2;
  wire       [253:0]  mdsMatrix_18_3;
  wire       [254:0]  mdsMatrix_18_4;
  wire       [254:0]  mdsMatrix_18_5;
  wire       [251:0]  mdsMatrix_18_6;
  wire       [251:0]  mdsMatrix_18_7;
  wire       [254:0]  mdsMatrix_18_8;
  wire       [254:0]  mdsMatrix_18_9;
  wire       [254:0]  mdsMatrix_18_10;
  wire       [254:0]  mdsMatrix_18_11;
  wire       [254:0]  mdsMatrix_19_0;
  wire       [254:0]  mdsMatrix_19_1;
  wire       [254:0]  mdsMatrix_19_2;
  wire       [254:0]  mdsMatrix_19_3;
  wire       [253:0]  mdsMatrix_19_4;
  wire       [251:0]  mdsMatrix_19_5;
  wire       [253:0]  mdsMatrix_19_6;
  wire       [254:0]  mdsMatrix_19_7;
  wire       [252:0]  mdsMatrix_19_8;
  wire       [253:0]  mdsMatrix_19_9;
  wire       [252:0]  mdsMatrix_19_10;
  wire       [254:0]  mdsMatrix_19_11;
  wire       [254:0]  mdsMatrix_20_0;
  wire       [254:0]  mdsMatrix_20_1;
  wire       [252:0]  mdsMatrix_20_2;
  wire       [253:0]  mdsMatrix_20_3;
  wire       [252:0]  mdsMatrix_20_4;
  wire       [253:0]  mdsMatrix_20_5;
  wire       [254:0]  mdsMatrix_20_6;
  wire       [252:0]  mdsMatrix_20_7;
  wire       [254:0]  mdsMatrix_20_8;
  wire       [251:0]  mdsMatrix_20_9;
  wire       [253:0]  mdsMatrix_20_10;
  wire       [252:0]  mdsMatrix_20_11;
  wire       [254:0]  mdsMatrix_21_0;
  wire       [254:0]  mdsMatrix_21_1;
  wire       [254:0]  mdsMatrix_21_2;
  wire       [254:0]  mdsMatrix_21_3;
  wire       [248:0]  mdsMatrix_21_4;
  wire       [254:0]  mdsMatrix_21_5;
  wire       [251:0]  mdsMatrix_21_6;
  wire       [254:0]  mdsMatrix_21_7;
  wire       [252:0]  mdsMatrix_21_8;
  wire       [254:0]  mdsMatrix_21_9;
  wire       [254:0]  mdsMatrix_21_10;
  wire       [253:0]  mdsMatrix_21_11;
  wire       [254:0]  mdsMatrix_22_0;
  wire       [254:0]  mdsMatrix_22_1;
  wire       [254:0]  mdsMatrix_22_2;
  wire       [254:0]  mdsMatrix_22_3;
  wire       [251:0]  mdsMatrix_22_4;
  wire       [252:0]  mdsMatrix_22_5;
  wire       [253:0]  mdsMatrix_22_6;
  wire       [253:0]  mdsMatrix_22_7;
  wire       [254:0]  mdsMatrix_22_8;
  wire       [253:0]  mdsMatrix_22_9;
  wire       [254:0]  mdsMatrix_22_10;
  wire       [254:0]  mdsMatrix_22_11;
  wire       [254:0]  mdsMatrix_23_0;
  wire       [250:0]  mdsMatrix_23_1;
  wire       [251:0]  mdsMatrix_23_2;
  wire       [252:0]  mdsMatrix_23_3;
  wire       [252:0]  mdsMatrix_23_4;
  wire       [252:0]  mdsMatrix_23_5;
  wire       [253:0]  mdsMatrix_23_6;
  wire       [253:0]  mdsMatrix_23_7;
  wire       [254:0]  mdsMatrix_23_8;
  wire       [254:0]  mdsMatrix_23_9;
  wire       [249:0]  mdsMatrix_23_10;
  wire       [253:0]  mdsMatrix_23_11;
  wire       [254:0]  mdsMatrix_24_0;
  wire       [253:0]  mdsMatrix_24_1;
  wire       [254:0]  mdsMatrix_24_2;
  wire       [253:0]  mdsMatrix_24_3;
  wire       [251:0]  mdsMatrix_24_4;
  wire       [254:0]  mdsMatrix_24_5;
  wire       [253:0]  mdsMatrix_24_6;
  wire       [253:0]  mdsMatrix_24_7;
  wire       [253:0]  mdsMatrix_24_8;
  wire       [253:0]  mdsMatrix_24_9;
  wire       [251:0]  mdsMatrix_24_10;
  wire       [253:0]  mdsMatrix_24_11;
  wire       [254:0]  mdsMatrix_25_0;
  wire       [254:0]  mdsMatrix_25_1;
  wire       [252:0]  mdsMatrix_25_2;
  wire       [250:0]  mdsMatrix_25_3;
  wire       [253:0]  mdsMatrix_25_4;
  wire       [252:0]  mdsMatrix_25_5;
  wire       [253:0]  mdsMatrix_25_6;
  wire       [253:0]  mdsMatrix_25_7;
  wire       [252:0]  mdsMatrix_25_8;
  wire       [253:0]  mdsMatrix_25_9;
  wire       [254:0]  mdsMatrix_25_10;
  wire       [254:0]  mdsMatrix_25_11;
  wire       [254:0]  mdsMatrix_26_0;
  wire       [253:0]  mdsMatrix_26_1;
  wire       [250:0]  mdsMatrix_26_2;
  wire       [250:0]  mdsMatrix_26_3;
  wire       [254:0]  mdsMatrix_26_4;
  wire       [253:0]  mdsMatrix_26_5;
  wire       [254:0]  mdsMatrix_26_6;
  wire       [252:0]  mdsMatrix_26_7;
  wire       [254:0]  mdsMatrix_26_8;
  wire       [251:0]  mdsMatrix_26_9;
  wire       [253:0]  mdsMatrix_26_10;
  wire       [253:0]  mdsMatrix_26_11;
  wire       [254:0]  mdsMatrix_27_0;
  wire       [254:0]  mdsMatrix_27_1;
  wire       [253:0]  mdsMatrix_27_2;
  wire       [253:0]  mdsMatrix_27_3;
  wire       [254:0]  mdsMatrix_27_4;
  wire       [253:0]  mdsMatrix_27_5;
  wire       [253:0]  mdsMatrix_27_6;
  wire       [254:0]  mdsMatrix_27_7;
  wire       [254:0]  mdsMatrix_27_8;
  wire       [252:0]  mdsMatrix_27_9;
  wire       [253:0]  mdsMatrix_27_10;
  wire       [252:0]  mdsMatrix_27_11;
  wire       [254:0]  mdsMatrix_28_0;
  wire       [251:0]  mdsMatrix_28_1;
  wire       [253:0]  mdsMatrix_28_2;
  wire       [254:0]  mdsMatrix_28_3;
  wire       [254:0]  mdsMatrix_28_4;
  wire       [250:0]  mdsMatrix_28_5;
  wire       [253:0]  mdsMatrix_28_6;
  wire       [254:0]  mdsMatrix_28_7;
  wire       [254:0]  mdsMatrix_28_8;
  wire       [254:0]  mdsMatrix_28_9;
  wire       [253:0]  mdsMatrix_28_10;
  wire       [253:0]  mdsMatrix_28_11;
  wire       [254:0]  mdsMatrix_29_0;
  wire       [254:0]  mdsMatrix_29_1;
  wire       [253:0]  mdsMatrix_29_2;
  wire       [254:0]  mdsMatrix_29_3;
  wire       [254:0]  mdsMatrix_29_4;
  wire       [253:0]  mdsMatrix_29_5;
  wire       [254:0]  mdsMatrix_29_6;
  wire       [254:0]  mdsMatrix_29_7;
  wire       [251:0]  mdsMatrix_29_8;
  wire       [253:0]  mdsMatrix_29_9;
  wire       [252:0]  mdsMatrix_29_10;
  wire       [253:0]  mdsMatrix_29_11;
  wire       [254:0]  mdsMatrix_30_0;
  wire       [253:0]  mdsMatrix_30_1;
  wire       [253:0]  mdsMatrix_30_2;
  wire       [249:0]  mdsMatrix_30_3;
  wire       [253:0]  mdsMatrix_30_4;
  wire       [254:0]  mdsMatrix_30_5;
  wire       [254:0]  mdsMatrix_30_6;
  wire       [254:0]  mdsMatrix_30_7;
  wire       [253:0]  mdsMatrix_30_8;
  wire       [254:0]  mdsMatrix_30_9;
  wire       [254:0]  mdsMatrix_30_10;
  wire       [252:0]  mdsMatrix_30_11;
  wire       [254:0]  mdsMatrix_31_0;
  wire       [252:0]  mdsMatrix_31_1;
  wire       [254:0]  mdsMatrix_31_2;
  wire       [253:0]  mdsMatrix_31_3;
  wire       [252:0]  mdsMatrix_31_4;
  wire       [254:0]  mdsMatrix_31_5;
  wire       [252:0]  mdsMatrix_31_6;
  wire       [254:0]  mdsMatrix_31_7;
  wire       [252:0]  mdsMatrix_31_8;
  wire       [253:0]  mdsMatrix_31_9;
  wire       [254:0]  mdsMatrix_31_10;
  wire       [254:0]  mdsMatrix_31_11;
  wire       [254:0]  mdsMatrix_32_0;
  wire       [254:0]  mdsMatrix_32_1;
  wire       [254:0]  mdsMatrix_32_2;
  wire       [254:0]  mdsMatrix_32_3;
  wire       [254:0]  mdsMatrix_32_4;
  wire       [251:0]  mdsMatrix_32_5;
  wire       [251:0]  mdsMatrix_32_6;
  wire       [253:0]  mdsMatrix_32_7;
  wire       [254:0]  mdsMatrix_32_8;
  wire       [254:0]  mdsMatrix_32_9;
  wire       [249:0]  mdsMatrix_32_10;
  wire       [252:0]  mdsMatrix_32_11;
  wire       [254:0]  mdsMatrix_33_0;
  wire       [254:0]  mdsMatrix_33_1;
  wire       [254:0]  mdsMatrix_33_2;
  wire       [253:0]  mdsMatrix_33_3;
  wire       [252:0]  mdsMatrix_33_4;
  wire       [254:0]  mdsMatrix_33_5;
  wire       [251:0]  mdsMatrix_33_6;
  wire       [252:0]  mdsMatrix_33_7;
  wire       [253:0]  mdsMatrix_33_8;
  wire       [251:0]  mdsMatrix_33_9;
  wire       [250:0]  mdsMatrix_33_10;
  wire       [251:0]  mdsMatrix_33_11;
  wire       [254:0]  mdsMatrix_34_0;
  wire       [253:0]  mdsMatrix_34_1;
  wire       [254:0]  mdsMatrix_34_2;
  wire       [252:0]  mdsMatrix_34_3;
  wire       [250:0]  mdsMatrix_34_4;
  wire       [254:0]  mdsMatrix_34_5;
  wire       [254:0]  mdsMatrix_34_6;
  wire       [254:0]  mdsMatrix_34_7;
  wire       [254:0]  mdsMatrix_34_8;
  wire       [253:0]  mdsMatrix_34_9;
  wire       [252:0]  mdsMatrix_34_10;
  wire       [254:0]  mdsMatrix_34_11;
  wire       [254:0]  mdsMatrix_35_0;
  wire       [253:0]  mdsMatrix_35_1;
  wire       [254:0]  mdsMatrix_35_2;
  wire       [254:0]  mdsMatrix_35_3;
  wire       [254:0]  mdsMatrix_35_4;
  wire       [252:0]  mdsMatrix_35_5;
  wire       [253:0]  mdsMatrix_35_6;
  wire       [253:0]  mdsMatrix_35_7;
  wire       [254:0]  mdsMatrix_35_8;
  wire       [252:0]  mdsMatrix_35_9;
  wire       [254:0]  mdsMatrix_35_10;
  wire       [254:0]  mdsMatrix_35_11;
  wire       [254:0]  mdsMatrix_36_0;
  wire       [254:0]  mdsMatrix_36_1;
  wire       [252:0]  mdsMatrix_36_2;
  wire       [248:0]  mdsMatrix_36_3;
  wire       [251:0]  mdsMatrix_36_4;
  wire       [254:0]  mdsMatrix_36_5;
  wire       [252:0]  mdsMatrix_36_6;
  wire       [253:0]  mdsMatrix_36_7;
  wire       [253:0]  mdsMatrix_36_8;
  wire       [253:0]  mdsMatrix_36_9;
  wire       [253:0]  mdsMatrix_36_10;
  wire       [253:0]  mdsMatrix_36_11;
  wire       [254:0]  mdsMatrix_37_0;
  wire       [251:0]  mdsMatrix_37_1;
  wire       [254:0]  mdsMatrix_37_2;
  wire       [254:0]  mdsMatrix_37_3;
  wire       [251:0]  mdsMatrix_37_4;
  wire       [253:0]  mdsMatrix_37_5;
  wire       [254:0]  mdsMatrix_37_6;
  wire       [254:0]  mdsMatrix_37_7;
  wire       [250:0]  mdsMatrix_37_8;
  wire       [254:0]  mdsMatrix_37_9;
  wire       [254:0]  mdsMatrix_37_10;
  wire       [253:0]  mdsMatrix_37_11;
  wire       [254:0]  mdsMatrix_38_0;
  wire       [253:0]  mdsMatrix_38_1;
  wire       [254:0]  mdsMatrix_38_2;
  wire       [253:0]  mdsMatrix_38_3;
  wire       [253:0]  mdsMatrix_38_4;
  wire       [254:0]  mdsMatrix_38_5;
  wire       [251:0]  mdsMatrix_38_6;
  wire       [253:0]  mdsMatrix_38_7;
  wire       [250:0]  mdsMatrix_38_8;
  wire       [254:0]  mdsMatrix_38_9;
  wire       [254:0]  mdsMatrix_38_10;
  wire       [254:0]  mdsMatrix_38_11;
  wire       [254:0]  mdsMatrix_39_0;
  wire       [254:0]  mdsMatrix_39_1;
  wire       [251:0]  mdsMatrix_39_2;
  wire       [249:0]  mdsMatrix_39_3;
  wire       [252:0]  mdsMatrix_39_4;
  wire       [252:0]  mdsMatrix_39_5;
  wire       [254:0]  mdsMatrix_39_6;
  wire       [253:0]  mdsMatrix_39_7;
  wire       [254:0]  mdsMatrix_39_8;
  wire       [254:0]  mdsMatrix_39_9;
  wire       [253:0]  mdsMatrix_39_10;
  wire       [254:0]  mdsMatrix_39_11;
  wire       [254:0]  mdsMatrix_40_0;
  wire       [254:0]  mdsMatrix_40_1;
  wire       [253:0]  mdsMatrix_40_2;
  wire       [254:0]  mdsMatrix_40_3;
  wire       [252:0]  mdsMatrix_40_4;
  wire       [254:0]  mdsMatrix_40_5;
  wire       [251:0]  mdsMatrix_40_6;
  wire       [254:0]  mdsMatrix_40_7;
  wire       [254:0]  mdsMatrix_40_8;
  wire       [253:0]  mdsMatrix_40_9;
  wire       [252:0]  mdsMatrix_40_10;
  wire       [250:0]  mdsMatrix_40_11;
  wire       [254:0]  mdsMatrix_41_0;
  wire       [254:0]  mdsMatrix_41_1;
  wire       [251:0]  mdsMatrix_41_2;
  wire       [254:0]  mdsMatrix_41_3;
  wire       [253:0]  mdsMatrix_41_4;
  wire       [254:0]  mdsMatrix_41_5;
  wire       [254:0]  mdsMatrix_41_6;
  wire       [254:0]  mdsMatrix_41_7;
  wire       [253:0]  mdsMatrix_41_8;
  wire       [253:0]  mdsMatrix_41_9;
  wire       [253:0]  mdsMatrix_41_10;
  wire       [253:0]  mdsMatrix_41_11;
  wire       [254:0]  mdsMatrix_42_0;
  wire       [252:0]  mdsMatrix_42_1;
  wire       [253:0]  mdsMatrix_42_2;
  wire       [250:0]  mdsMatrix_42_3;
  wire       [252:0]  mdsMatrix_42_4;
  wire       [253:0]  mdsMatrix_42_5;
  wire       [249:0]  mdsMatrix_42_6;
  wire       [254:0]  mdsMatrix_42_7;
  wire       [254:0]  mdsMatrix_42_8;
  wire       [253:0]  mdsMatrix_42_9;
  wire       [252:0]  mdsMatrix_42_10;
  wire       [254:0]  mdsMatrix_42_11;
  wire       [254:0]  mdsMatrix_43_0;
  wire       [252:0]  mdsMatrix_43_1;
  wire       [250:0]  mdsMatrix_43_2;
  wire       [254:0]  mdsMatrix_43_3;
  wire       [254:0]  mdsMatrix_43_4;
  wire       [254:0]  mdsMatrix_43_5;
  wire       [254:0]  mdsMatrix_43_6;
  wire       [253:0]  mdsMatrix_43_7;
  wire       [253:0]  mdsMatrix_43_8;
  wire       [249:0]  mdsMatrix_43_9;
  wire       [251:0]  mdsMatrix_43_10;
  wire       [254:0]  mdsMatrix_43_11;
  wire       [254:0]  mdsMatrix_44_0;
  wire       [254:0]  mdsMatrix_44_1;
  wire       [251:0]  mdsMatrix_44_2;
  wire       [253:0]  mdsMatrix_44_3;
  wire       [253:0]  mdsMatrix_44_4;
  wire       [252:0]  mdsMatrix_44_5;
  wire       [251:0]  mdsMatrix_44_6;
  wire       [254:0]  mdsMatrix_44_7;
  wire       [253:0]  mdsMatrix_44_8;
  wire       [253:0]  mdsMatrix_44_9;
  wire       [254:0]  mdsMatrix_44_10;
  wire       [252:0]  mdsMatrix_44_11;
  wire       [254:0]  mdsMatrix_45_0;
  wire       [254:0]  mdsMatrix_45_1;
  wire       [254:0]  mdsMatrix_45_2;
  wire       [254:0]  mdsMatrix_45_3;
  wire       [254:0]  mdsMatrix_45_4;
  wire       [253:0]  mdsMatrix_45_5;
  wire       [253:0]  mdsMatrix_45_6;
  wire       [254:0]  mdsMatrix_45_7;
  wire       [252:0]  mdsMatrix_45_8;
  wire       [249:0]  mdsMatrix_45_9;
  wire       [254:0]  mdsMatrix_45_10;
  wire       [254:0]  mdsMatrix_45_11;
  wire       [254:0]  mdsMatrix_46_0;
  wire       [253:0]  mdsMatrix_46_1;
  wire       [252:0]  mdsMatrix_46_2;
  wire       [254:0]  mdsMatrix_46_3;
  wire       [253:0]  mdsMatrix_46_4;
  wire       [254:0]  mdsMatrix_46_5;
  wire       [254:0]  mdsMatrix_46_6;
  wire       [254:0]  mdsMatrix_46_7;
  wire       [254:0]  mdsMatrix_46_8;
  wire       [254:0]  mdsMatrix_46_9;
  wire       [252:0]  mdsMatrix_46_10;
  wire       [253:0]  mdsMatrix_46_11;
  wire       [254:0]  mdsMatrix_47_0;
  wire       [251:0]  mdsMatrix_47_1;
  wire       [249:0]  mdsMatrix_47_2;
  wire       [254:0]  mdsMatrix_47_3;
  wire       [251:0]  mdsMatrix_47_4;
  wire       [253:0]  mdsMatrix_47_5;
  wire       [254:0]  mdsMatrix_47_6;
  wire       [254:0]  mdsMatrix_47_7;
  wire       [254:0]  mdsMatrix_47_8;
  wire       [253:0]  mdsMatrix_47_9;
  wire       [254:0]  mdsMatrix_47_10;
  wire       [254:0]  mdsMatrix_47_11;
  wire       [254:0]  mdsMatrix_48_0;
  wire       [251:0]  mdsMatrix_48_1;
  wire       [253:0]  mdsMatrix_48_2;
  wire       [254:0]  mdsMatrix_48_3;
  wire       [253:0]  mdsMatrix_48_4;
  wire       [253:0]  mdsMatrix_48_5;
  wire       [254:0]  mdsMatrix_48_6;
  wire       [252:0]  mdsMatrix_48_7;
  wire       [253:0]  mdsMatrix_48_8;
  wire       [253:0]  mdsMatrix_48_9;
  wire       [254:0]  mdsMatrix_48_10;
  wire       [254:0]  mdsMatrix_48_11;
  wire       [254:0]  mdsMatrix_49_0;
  wire       [251:0]  mdsMatrix_49_1;
  wire       [254:0]  mdsMatrix_49_2;
  wire       [254:0]  mdsMatrix_49_3;
  wire       [253:0]  mdsMatrix_49_4;
  wire       [254:0]  mdsMatrix_49_5;
  wire       [252:0]  mdsMatrix_49_6;
  wire       [254:0]  mdsMatrix_49_7;
  wire       [252:0]  mdsMatrix_49_8;
  wire       [254:0]  mdsMatrix_49_9;
  wire       [253:0]  mdsMatrix_49_10;
  wire       [254:0]  mdsMatrix_49_11;
  wire       [254:0]  mdsMatrix_50_0;
  wire       [251:0]  mdsMatrix_50_1;
  wire       [254:0]  mdsMatrix_50_2;
  wire       [254:0]  mdsMatrix_50_3;
  wire       [252:0]  mdsMatrix_50_4;
  wire       [253:0]  mdsMatrix_50_5;
  wire       [253:0]  mdsMatrix_50_6;
  wire       [252:0]  mdsMatrix_50_7;
  wire       [254:0]  mdsMatrix_50_8;
  wire       [254:0]  mdsMatrix_50_9;
  wire       [252:0]  mdsMatrix_50_10;
  wire       [252:0]  mdsMatrix_50_11;
  wire       [254:0]  mdsMatrix_51_0;
  wire       [254:0]  mdsMatrix_51_1;
  wire       [253:0]  mdsMatrix_51_2;
  wire       [254:0]  mdsMatrix_51_3;
  wire       [252:0]  mdsMatrix_51_4;
  wire       [254:0]  mdsMatrix_51_5;
  wire       [253:0]  mdsMatrix_51_6;
  wire       [254:0]  mdsMatrix_51_7;
  wire       [252:0]  mdsMatrix_51_8;
  wire       [253:0]  mdsMatrix_51_9;
  wire       [254:0]  mdsMatrix_51_10;
  wire       [254:0]  mdsMatrix_51_11;
  wire       [254:0]  mdsMatrix_52_0;
  wire       [254:0]  mdsMatrix_52_1;
  wire       [253:0]  mdsMatrix_52_2;
  wire       [252:0]  mdsMatrix_52_3;
  wire       [253:0]  mdsMatrix_52_4;
  wire       [253:0]  mdsMatrix_52_5;
  wire       [253:0]  mdsMatrix_52_6;
  wire       [253:0]  mdsMatrix_52_7;
  wire       [254:0]  mdsMatrix_52_8;
  wire       [254:0]  mdsMatrix_52_9;
  wire       [252:0]  mdsMatrix_52_10;
  wire       [254:0]  mdsMatrix_52_11;
  wire       [254:0]  mdsMatrix_53_0;
  wire       [250:0]  mdsMatrix_53_1;
  wire       [253:0]  mdsMatrix_53_2;
  wire       [254:0]  mdsMatrix_53_3;
  wire       [251:0]  mdsMatrix_53_4;
  wire       [254:0]  mdsMatrix_53_5;
  wire       [253:0]  mdsMatrix_53_6;
  wire       [254:0]  mdsMatrix_53_7;
  wire       [254:0]  mdsMatrix_53_8;
  wire       [254:0]  mdsMatrix_53_9;
  wire       [252:0]  mdsMatrix_53_10;
  wire       [254:0]  mdsMatrix_53_11;
  wire       [254:0]  mdsMatrix_54_0;
  wire       [254:0]  mdsMatrix_54_1;
  wire       [253:0]  mdsMatrix_54_2;
  wire       [254:0]  mdsMatrix_54_3;
  wire       [254:0]  mdsMatrix_54_4;
  wire       [254:0]  mdsMatrix_54_5;
  wire       [253:0]  mdsMatrix_54_6;
  wire       [253:0]  mdsMatrix_54_7;
  wire       [252:0]  mdsMatrix_54_8;
  wire       [253:0]  mdsMatrix_54_9;
  wire       [253:0]  mdsMatrix_54_10;
  wire       [254:0]  mdsMatrix_54_11;
  wire       [254:0]  mdsMatrix_55_0;
  wire       [253:0]  mdsMatrix_55_1;
  wire       [254:0]  mdsMatrix_55_2;
  wire       [254:0]  mdsMatrix_55_3;
  wire       [254:0]  mdsMatrix_55_4;
  wire       [252:0]  mdsMatrix_55_5;
  wire       [253:0]  mdsMatrix_55_6;
  wire       [246:0]  mdsMatrix_55_7;
  wire       [252:0]  mdsMatrix_55_8;
  wire       [254:0]  mdsMatrix_55_9;
  wire       [253:0]  mdsMatrix_55_10;
  wire       [251:0]  mdsMatrix_55_11;
  wire       [254:0]  mdsMatrix_56_0;
  wire       [254:0]  mdsMatrix_56_1;
  wire       [254:0]  mdsMatrix_56_2;
  wire       [253:0]  mdsMatrix_56_3;
  wire       [253:0]  mdsMatrix_56_4;
  wire       [249:0]  mdsMatrix_56_5;
  wire       [253:0]  mdsMatrix_56_6;
  wire       [254:0]  mdsMatrix_56_7;
  wire       [254:0]  mdsMatrix_56_8;
  wire       [252:0]  mdsMatrix_56_9;
  wire       [254:0]  mdsMatrix_56_10;
  wire       [247:0]  mdsMatrix_56_11;
  wire       [5:0]    tempAddrVec_0;
  wire       [5:0]    tempAddrVec_1;
  wire       [5:0]    tempAddrVec_2;
  wire       [5:0]    tempAddrVec_3;
  wire       [5:0]    tempAddrVec_4;
  wire       [5:0]    tempAddrVec_5;
  wire       [5:0]    tempAddrVec_6;
  wire       [5:0]    tempAddrVec_7;
  wire       [5:0]    tempAddrVec_8;
  wire       [5:0]    tempAddrVec_9;
  wire       [5:0]    tempAddrVec_10;
  wire       [5:0]    tempAddrVec_11;
  reg        [5:0]    io_addr_regNext;
  reg        [5:0]    io_addr_regNext_1;
  reg        [5:0]    io_addr_regNext_2;
  reg        [5:0]    io_addr_regNext_3;
  reg        [5:0]    io_addr_regNext_4;
  reg        [5:0]    io_addr_regNext_5;
  reg        [5:0]    io_addr_regNext_6;
  reg        [5:0]    io_addr_regNext_7;
  reg        [5:0]    io_addr_regNext_8;
  reg        [5:0]    io_addr_regNext_9;
  reg        [5:0]    io_addr_regNext_10;
  reg        [5:0]    io_addr_regNext_11;
  reg [254:0] mdsMem_0 [0:56];
  reg [254:0] mdsMem_1 [0:56];
  reg [254:0] mdsMem_2 [0:56];
  reg [254:0] mdsMem_3 [0:56];
  reg [254:0] mdsMem_4 [0:56];
  reg [254:0] mdsMem_5 [0:56];
  reg [254:0] mdsMem_6 [0:56];
  reg [254:0] mdsMem_7 [0:56];
  reg [254:0] mdsMem_8 [0:56];
  reg [254:0] mdsMem_9 [0:56];
  reg [254:0] mdsMem_10 [0:56];
  reg [254:0] mdsMem_11 [0:56];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  assign _zz_io_data_5 = 1'b1;
  assign _zz_io_data_6 = 1'b1;
  assign _zz_io_data_7 = 1'b1;
  assign _zz_io_data_8 = 1'b1;
  assign _zz_io_data_9 = 1'b1;
  assign _zz_io_data_10 = 1'b1;
  assign _zz_io_data_11 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_5.bin",mdsMem_5);
  end
  always @(posedge clk) begin
    if(_zz_io_data_5) begin
      _zz_mdsMem_5_port0 <= mdsMem_5[tempAddrVec_5];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_6.bin",mdsMem_6);
  end
  always @(posedge clk) begin
    if(_zz_io_data_6) begin
      _zz_mdsMem_6_port0 <= mdsMem_6[tempAddrVec_6];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_7.bin",mdsMem_7);
  end
  always @(posedge clk) begin
    if(_zz_io_data_7) begin
      _zz_mdsMem_7_port0 <= mdsMem_7[tempAddrVec_7];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_8.bin",mdsMem_8);
  end
  always @(posedge clk) begin
    if(_zz_io_data_8) begin
      _zz_mdsMem_8_port0 <= mdsMem_8[tempAddrVec_8];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_9.bin",mdsMem_9);
  end
  always @(posedge clk) begin
    if(_zz_io_data_9) begin
      _zz_mdsMem_9_port0 <= mdsMem_9[tempAddrVec_9];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_10.bin",mdsMem_10);
  end
  always @(posedge clk) begin
    if(_zz_io_data_10) begin
      _zz_mdsMem_10_port0 <= mdsMem_10[tempAddrVec_10];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_27_mdsMem_11.bin",mdsMem_11);
  end
  always @(posedge clk) begin
    if(_zz_io_data_11) begin
      _zz_mdsMem_11_port0 <= mdsMem_11[tempAddrVec_11];
    end
  end

  assign mdsMatrix_0_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_0_1 = 255'h42047a37f7b388d1d8d435acc93ef61907614c5062735834822d956b2e486795;
  assign mdsMatrix_0_2 = 255'h55a94a22b3ed12486a4ff36778c9dd4978fa2c8b0db48fa402a5f58531f4fa74;
  assign mdsMatrix_0_3 = 254'h29daa09e4dc602187e687e401b0133efd1218025953188144af7629ca239a9ed;
  assign mdsMatrix_0_4 = 254'h31a8532d2e9885b139a50efda7b69b0a012d6c6b18e3d8f07f1b78bab5cf47e4;
  assign mdsMatrix_0_5 = 254'h2278e5c54cfdcc1d235d47c7f3f2813c21bb8329c88e28432f6d5b45080e246b;
  assign mdsMatrix_0_6 = 252'hfee22e77489943b6575f84a0b9ae2b9eddb4c1987277431f4bd11b54fa44e49;
  assign mdsMatrix_0_7 = 255'h631869cb5ff08a44ef9e6af537cf976a12e35eec0859b09efe8f3a529019e863;
  assign mdsMatrix_0_8 = 255'h68533d03208d580f068d1890bbc9a4d5adddc3dbf22f06119bcdda5515a4b85a;
  assign mdsMatrix_0_9 = 253'h1e59787b25d0399007a3913331a28ab9a9a4123af917c19dd66deab1ae612f27;
  assign mdsMatrix_0_10 = 254'h2b1310fc9c7b2e5de571eeeb9b2be654c70ff72963a29c8161cb5dc5da674abe;
  assign mdsMatrix_0_11 = 254'h2de89631a8b9b66cb00ec7169e898514bf95f76705de03973a54b1dc8c4840f5;
  assign mdsMatrix_1_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_1_1 = 254'h2c7b92479337cc847a55896681ed519aff8229d640f3d9605988e5fab71d837a;
  assign mdsMatrix_1_2 = 255'h49a274feac48d3607d14aca83390470862635e29afa9e29033ebbd3eb3edf1b8;
  assign mdsMatrix_1_3 = 255'h4cddcfdeb66d74557ab905757e2a14cafc838546685ed9ae80feeec0215922a6;
  assign mdsMatrix_1_4 = 251'h48b0dfe7dca6939ff4c40b203e1dd4ec7e51ecd87a7b47a2a160f296cb10bac;
  assign mdsMatrix_1_5 = 255'h4d2b461de9852f2424c69a8914560b8e4d75fb672ec71df9bb0face3ad005a35;
  assign mdsMatrix_1_6 = 255'h44236035c883d40426fc65636da9dee2c68a59de05dffef51cf2a2eb25191c9e;
  assign mdsMatrix_1_7 = 253'h10e84c53cb4ad5fe49def19b8b0bbed851e96a36ce1d9c79d7f7dc75fd3aaeb1;
  assign mdsMatrix_1_8 = 255'h647cd4f3bf3aecc587278b77adaa6bbf13807bba6d4c3d217ad8d2b897fbd75b;
  assign mdsMatrix_1_9 = 255'h5b8bccb0df83be11136c56b792be72a9333c66e8e5b762af11f6c62d0a3674ee;
  assign mdsMatrix_1_10 = 250'h26c8261a3763c640a6bac580b4dc7db7b943bd02dbe5a6ca5af77e2ebb08736;
  assign mdsMatrix_1_11 = 253'h10d6c2685ee3f1c276322e3ea7df5d919d166f8cb032584c99f0a9fead9a4a2c;
  assign mdsMatrix_2_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_2_1 = 253'h1e28fa627efdff879196591413e1e33ecfba0d7a34aae3dd0cd5342b75822122;
  assign mdsMatrix_2_2 = 254'h2e4a0f7df9bb02bf2e52c6f916639bb1557a1be044c03827d0d64f1f2d589b5e;
  assign mdsMatrix_2_3 = 254'h281dfac2bb025af4930d641092c47d5eb3d0b9d2cd3420b12ca395bbaeef705b;
  assign mdsMatrix_2_4 = 254'h3a65119082fb6604996afc1b8e78e599dd951f92b2329ed5c482548175b819b9;
  assign mdsMatrix_2_5 = 253'h1a9eaeb793e51773e681abe627b2fa425d62c2a5ce9d79f06f420ae900b75211;
  assign mdsMatrix_2_6 = 255'h497b7e435f7890df5c3d7a2d8a9943dfdfd6a17a1df09f7885efb407e89ee850;
  assign mdsMatrix_2_7 = 253'h1e4c55ea120e6ec18cf651cd9702cf75c130e652e42ed97bef41d93316e75e87;
  assign mdsMatrix_2_8 = 252'hb4105059d94821158b7e8f61ef4ea5e19ee6515aeabb34351d9957034d35ab0;
  assign mdsMatrix_2_9 = 250'h32a651b36979ee2460ce122ee77ea71681336ef03f669bcfeb9151a1c7c6acc;
  assign mdsMatrix_2_10 = 252'he2e250e8312856e3e5d34ed4eadd9f37f3d6e27f9844143ea4d28c3c3794fe7;
  assign mdsMatrix_2_11 = 255'h6fafeb1bf3cb52cf80c0b8add9ce9d6afa92a77f0a61acac240124f929f7e67b;
  assign mdsMatrix_3_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_3_1 = 253'h10a758565e899a7ecd7e1c48d3688a73d68ee67632738085ebc22fd85542a8d9;
  assign mdsMatrix_3_2 = 254'h2126576370dd0094d7f69bac3332af9462dfc089b9c29edc60672d7e2152daad;
  assign mdsMatrix_3_3 = 255'h41a0da384c46e7c55faad1840b8bc1fe79d67877fffa7751743e8d68bd997fc2;
  assign mdsMatrix_3_4 = 255'h67c6235b58d29c87d6c563e4ddf67091d6662fe07820834f979fbcecb5eed8a1;
  assign mdsMatrix_3_5 = 254'h2dacfaf7ccc49e47fe534ce800be8c7a79044b771f623a2ae4d0f21f4936a0f1;
  assign mdsMatrix_3_6 = 254'h39882a8dd537475a9a1598ab262da7db01d38bbebb496a6bfee7b6bc284e9316;
  assign mdsMatrix_3_7 = 252'h87aa1082391c70e219ee9f3777081e95105d8b12ba673f5e1e59e1183c1a37a;
  assign mdsMatrix_3_8 = 254'h26f5831d95037a5c76f053a3fc1169cdb074ae37a697a1140010a2382de1a978;
  assign mdsMatrix_3_9 = 255'h4d638416e7012ed16a8a961c98d40a4e0555102b8a01e30622033bc933f557ac;
  assign mdsMatrix_3_10 = 255'h720e2c7710a327051c6edfd19d9ac222025bf2bc83421e6dbfdb512fef9e854d;
  assign mdsMatrix_3_11 = 255'h73bf1906474640432d92a600dd20bdff5c098e6136a61d953810c071fc197da6;
  assign mdsMatrix_4_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_4_1 = 253'h1ce47670f185bfb4cdb71390c722ba2a3bc07cdf3afb852842f6747fe10c6d44;
  assign mdsMatrix_4_2 = 255'h556981491e35af7440acde2f33b3fa71e81899d76a898ad2f84e1c75f8aa4449;
  assign mdsMatrix_4_3 = 253'h125d9d7a240a6e4426f84d8f91e1952d5f55a713382fd412237d94f7d05dbd3c;
  assign mdsMatrix_4_4 = 254'h36a8d61ee9facd49f400754b07dc05f9aaaf4d11ad2783375ae7d56bd3a173e0;
  assign mdsMatrix_4_5 = 252'hab005f55f66213624536968a59d9a570979e8dae1d9c34434024c321c5ee8fa;
  assign mdsMatrix_4_6 = 253'h113ff1d91bdd9d9f6cce1321bb9f167b55995f8d4d7ebc77aceedc37378927e3;
  assign mdsMatrix_4_7 = 255'h73cd5094e5395cc4fd3bfdd71ad893f471ad4ea5ffc65b266c0d8d43c4d04799;
  assign mdsMatrix_4_8 = 255'h4654dab818d24828410645480de37138c72e06b017331a0c73689a5b6d107bd7;
  assign mdsMatrix_4_9 = 253'h1c0442f99174f5e6386a2fa47190c762c3d4be5d844dcdc1d102ab8132e7120c;
  assign mdsMatrix_4_10 = 252'h87220509ad14c33d306e75b1d62491088ed9700f22aa40960ae81704766111f;
  assign mdsMatrix_4_11 = 255'h5fd44a4f479cf95aaeede27630bce564c010715f3890d157118396eb91996058;
  assign mdsMatrix_5_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_5_1 = 255'h6bab001744a92a11baccd784bee4bba8c2a7680d88a3dc37739ef9eee18fa6f5;
  assign mdsMatrix_5_2 = 255'h56cab18244f554205b5d18b1b83fba5cb6dfc179797c2ab759a052f88d2bbe5f;
  assign mdsMatrix_5_3 = 254'h235764cddbd31656e298290ea1c46d43b1c3cb938927b202df1c170d09edff08;
  assign mdsMatrix_5_4 = 253'h18170fe136bf10f059addf265745f2d926c896cb65a70544ce0d3e58cf8ddaab;
  assign mdsMatrix_5_5 = 255'h68440cdd000fded848d22bd4d83df4648c4123df575451b5c5ee2f61c7ee0517;
  assign mdsMatrix_5_6 = 252'hd5c881138b6ace390dac403eb9cdfdf727056fa6068bde0f62fac710c2322b4;
  assign mdsMatrix_5_7 = 250'h2998c2275fd4d36b3f6da9d790451169c28fdb2b222613db83a1c5d948967c7;
  assign mdsMatrix_5_8 = 248'ha3eb5eb9b69fb4d25d954dd42ba89fb0cad6d1bef04b4b25d35bf2646c0551;
  assign mdsMatrix_5_9 = 254'h3089baf441bcb66d5314ddb0c63fc0b2d04e2d37a72432d3a9417d00bbb5643f;
  assign mdsMatrix_5_10 = 255'h68149eae6e2b56a8aa9505e47ab468063006b9b887df0ff4fd00129ae3e895fb;
  assign mdsMatrix_5_11 = 254'h32bcb103d5758e1723f516dbe09e5c7c15c69a8006c9f87fc0a4b6dcb3acf46e;
  assign mdsMatrix_6_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_6_1 = 255'h6485aae68ddc31cb1de9e1569fe24ebb501bf9696832a548f6412f44d97bb8fd;
  assign mdsMatrix_6_2 = 252'hc4f7ed87d391011c857042d6221a5ddeedabdb4ab04799e1ecdcbf0972edb35;
  assign mdsMatrix_6_3 = 254'h23da21d0bef1487c03fd80ba16f790327484883a7df71ce84ce3d81538292a0c;
  assign mdsMatrix_6_4 = 255'h6f191e17721caae52a66b0ada7b8c7b88af78120f4224c1ac2d503a5bf552a5f;
  assign mdsMatrix_6_5 = 253'h1bca9ac9b2fd982046982dec2fd719555f5159de4c8d3fba2ffef48bbb94fa06;
  assign mdsMatrix_6_6 = 254'h222877a0a4b4df25d4946952567b6e94d09e64472428b0545f18965fedd4a299;
  assign mdsMatrix_6_7 = 250'h3d5ce9177109f3c6be138ed5df70f484e1e65b088f609efd8c64deedf1c9eef;
  assign mdsMatrix_6_8 = 255'h6ae5f1ea670e5323457c78c957aa7d9457665448ab64b05476a632ae491c097d;
  assign mdsMatrix_6_9 = 252'hf18ac9e1dc1852107d6880d05dda4f89e05d6a02c51e45feafd4593a3055139;
  assign mdsMatrix_6_10 = 251'h4bd1248f2983c244d6c65be01254a3798570b911d9dbed102165ec507f2fc4d;
  assign mdsMatrix_6_11 = 254'h256863cc559dc44c17a2c8db1cfbdf063fdc8b6216fa1e30f52fcc5b79407648;
  assign mdsMatrix_7_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_7_1 = 253'h18e711db5bb3567d66eb14fdf2818ebba89fb7a88dbde0bb5fefa65387e3fc41;
  assign mdsMatrix_7_2 = 254'h2806178350ae91c3afa702364d84325ae2b8616b0512caadffb3612de0ea77b5;
  assign mdsMatrix_7_3 = 254'h24d8f3047cc6c887eb6eac9e3895932785d34af5c6d47f0bc32f4766e5d379e5;
  assign mdsMatrix_7_4 = 255'h67e46849c4a4e5dcdec658a10d37688b27c770defc0468c0346f1b37d155996d;
  assign mdsMatrix_7_5 = 254'h2c1441c4b8a061f4dbdea6e796c10793295fa6d4f3a7a9b7a06a022c1687ef52;
  assign mdsMatrix_7_6 = 254'h22f5607177e20953cfefd2210cf4f86d20c4a7b85f846ac182d14b7350e8c5a8;
  assign mdsMatrix_7_7 = 255'h5febe99b92d349b42b436f028f1237856582bce085f4a8e019f78a56e130dd1b;
  assign mdsMatrix_7_8 = 255'h50ca10f0ccb8c869b6dc03db91796fd86efdb6c3f0c81637e069ae08f8e1870e;
  assign mdsMatrix_7_9 = 254'h27d71f821ac0f855ad02cefdc50791dfd1a29e66543384a4f15b259b7b8faffa;
  assign mdsMatrix_7_10 = 254'h2b90d5f88d17359e4175fa305f29a896dff512352da336118467ff4312c8f383;
  assign mdsMatrix_7_11 = 254'h20097915285ff6eef29eed3ae5a8e275078b0a1ec4c1d9582aecfe5f38accf0c;
  assign mdsMatrix_8_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_8_1 = 255'h5df4763e6c37ea2395314039fdb4ab0c99fe24cf82fa15fffc86a3a4629d840e;
  assign mdsMatrix_8_2 = 255'h4bd821842f5490783488b2396a28736ffdb32939f6506696641e5535f63b234a;
  assign mdsMatrix_8_3 = 255'h619beb865bd5d1dace5abdb27333c2957847ba165c9e28ccd84da190838c03fd;
  assign mdsMatrix_8_4 = 254'h30477dc313dc4aaa532a6e2609418f024f412b9e091787ab7ad8049971daa7fb;
  assign mdsMatrix_8_5 = 255'h476b67d964bcfa69e21f2947ed779069066b48e9c59a9a12814750424dc73b50;
  assign mdsMatrix_8_6 = 255'h42886ed2091b67a3bd90fa4595e10cca39a12c8b291e8686ac2a5c95bc7070c2;
  assign mdsMatrix_8_7 = 249'h1ae42e0e7ee1a0b17e436dc8f49e6c0b378373e4686ad9c87bdfd425b436681;
  assign mdsMatrix_8_8 = 253'h10462e2f82528d06d0a4cbe8daf52daa30c3dc1f198afc3bacd8dc629637860a;
  assign mdsMatrix_8_9 = 252'hac8dc8382cc3c34d0984e0286cfd12bd61f0c2fe4758ccf142f308095a4db4c;
  assign mdsMatrix_8_10 = 254'h2932aa33ee181c81a38c2782f8fc06404201c921577366eff15b0be3db015c80;
  assign mdsMatrix_8_11 = 254'h262add18d12592ba6a7e3074ade3d05d9b52699c9cd5f57e61d49aba141319a0;
  assign mdsMatrix_9_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_9_1 = 253'h11601fbc144cacd1e7de40d3995dca16fbd7fbdbba45c500e9ff69697fb82295;
  assign mdsMatrix_9_2 = 254'h378726ef7423676f549198a4dd575aae127734ff4a1039bb9b1abbb640d94fc6;
  assign mdsMatrix_9_3 = 255'h63d5b3b25fc3fccd70b27834e8a6900f67cac74601e7793316258386af32a9af;
  assign mdsMatrix_9_4 = 254'h266dd7ccdd9bdd823aab181e53241dc295b1ca08099866c2fc43b659df7455a4;
  assign mdsMatrix_9_5 = 253'h18cface6efe8133099d303ff38e8c8eb58249ec8ce8a346326fd0ef738720345;
  assign mdsMatrix_9_6 = 255'h723d4c7e56b4e458a9ff8b400f41319bae60e0b1a70bde18582f4e8dee0447a9;
  assign mdsMatrix_9_7 = 254'h35ef85f610402d9991c6a8bca62264122a33a9211432ce686e2ef538e6f356d5;
  assign mdsMatrix_9_8 = 253'h137058fe794d2ff4a1864d7017eef03c9f42290a3f7bafeb7ea31ae51d31c9ea;
  assign mdsMatrix_9_9 = 253'h1d82928e118b74b1315bbae1713c1f7a84078c3fac9399ffa43d17d13e7c32a1;
  assign mdsMatrix_9_10 = 254'h33ca93c21c716f85ad4bb910a8beeb61b73e3ccb95fea3b0a3b5ac41af46b97f;
  assign mdsMatrix_9_11 = 255'h59c403b77ce3cc91e4975238347e7f19f04b9679fddd713a1254c4677f409448;
  assign mdsMatrix_10_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_10_1 = 255'h42160d27cdff9f24a1c4f664c22686ba00823b5a3aa631e692ad3c9e9acc6110;
  assign mdsMatrix_10_2 = 255'h607a6e92ec439cae8541fbb4498c0cce2b623657aea87d4c0b7100cf2d412507;
  assign mdsMatrix_10_3 = 255'h6a54f1b17fb7ed329860f7e4149d40ed4f1b19c2ef49a3956aee8f02f95d29c4;
  assign mdsMatrix_10_4 = 252'h9fda2f0770731d55000235b2f97a89fb444a94416038aaa045c499c99b9d3e4;
  assign mdsMatrix_10_5 = 255'h41a120b5d1eb7547e61b7e90f5dae458e03c810546e387b83d3843d72680e56e;
  assign mdsMatrix_10_6 = 253'h1a28231bb3f7c470dd4ba8988b290b43bc5692a1ee1918ff7c85d8c63a6a92d8;
  assign mdsMatrix_10_7 = 254'h3218131c435c54c72920b355d2d2d3d60398a05c421b6967ecc36de9347edcaf;
  assign mdsMatrix_10_8 = 255'h6d1a87064b0fe88656974db47c6cbf2d7ed4c4d394b702c75fd11c434441ccde;
  assign mdsMatrix_10_9 = 254'h2a62f184a40000fc4f982cdbd5b4d9d5da47843030f98713d41fe15e6c7743e1;
  assign mdsMatrix_10_10 = 253'h117158f5bab34db91e457772418f9f7738f735395ff55a3b08332efd85538feb;
  assign mdsMatrix_10_11 = 255'h5864fd00d39db39bda835d29bf09500f429ddc15695cfa9dcc9908b0a3a05dd9;
  assign mdsMatrix_11_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_11_1 = 254'h2505560f72198d31161497c5b843f20441cc330fd67173a694e8b1728198dafc;
  assign mdsMatrix_11_2 = 252'hcf31a662af0218bb9ebce259079a79bba540c9971fe1ff48b4cdb8916dcc5d4;
  assign mdsMatrix_11_3 = 255'h54349a10c7583181e73af88e88b17ad6fa4a8d9405514b36c5aae1edf52827dc;
  assign mdsMatrix_11_4 = 255'h48513c65adfb49bc3ab36189f4b2636a734b9ff154436b02e9a4b1974dc76649;
  assign mdsMatrix_11_5 = 255'h512c8a1aeaf73ea581b9cd4090101fe00cefdb676aeb0c4dc3791479e5641e6b;
  assign mdsMatrix_11_6 = 253'h1cbcb6039be1dc584dfdd29ea46be9c4e08d51b8328956b7948409b214478cb8;
  assign mdsMatrix_11_7 = 255'h60437466d9310d081debca7bb1faa1b17aba281c95942138a5469ce797e4c713;
  assign mdsMatrix_11_8 = 253'h1db128eb3eef92ba87517f8d60f3bdc84a023a7e50583872025d8380181ba04a;
  assign mdsMatrix_11_9 = 253'h170442d9d076f9a5e1782010393aedbcbde3bcabe6904674e0c0e3881d108eff;
  assign mdsMatrix_11_10 = 254'h21aaad49095121b15e071f061dd8e18295b2afb367810dd14cf285bdd6212be0;
  assign mdsMatrix_11_11 = 254'h245ce5c005296083510988e98159357a69913be2e6a3910fba372f2a5488eee7;
  assign mdsMatrix_12_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_12_1 = 255'h41ded6716a174c5681ee6c88cd8a6aaa00ec37a6d24e70f27255e93979edde55;
  assign mdsMatrix_12_2 = 255'h5cfe7283172d1fdb8c80dac070a86415f1ae38f076aa1ee48a76a6aed67025f5;
  assign mdsMatrix_12_3 = 255'h46e7b1301e0c9d95f210093925b257ce4d7caf1b3e1a0b3595fcfcaaab715a8d;
  assign mdsMatrix_12_4 = 253'h19765d63caaa73a41cd5ec9b249d0470127a7b403f07bf3c25082d5ca8419ab8;
  assign mdsMatrix_12_5 = 254'h37459a7bd14b199dfcc24bb97156a77b0f2d68e8d3d7bfafbe086cf95230ba8b;
  assign mdsMatrix_12_6 = 255'h58797b19ab9f84e73f7edf64cbcceecd4065e1e81400b7b59b8dafaf2ca03c7e;
  assign mdsMatrix_12_7 = 254'h2c4f3f4c75bf082f9f0b49d473f8a7072b22431bef5920a4ee432d9e3ad52d5a;
  assign mdsMatrix_12_8 = 255'h43bc5964c510e58237fb38f1efdd11e74292a07c2220e47d0340c05f82e677f5;
  assign mdsMatrix_12_9 = 253'h106abd23f4dc5772f9b8917d37b1b6eeca272d3cd51fd6a344ce2db8d554cfc0;
  assign mdsMatrix_12_10 = 255'h682fcdf41011afac1196c64d0120525b81eb698444553487761a8f1c35286b48;
  assign mdsMatrix_12_11 = 255'h6e0119a8f68a4457b012c2f78253ca9dcebc82a627802f35576900307a0753bb;
  assign mdsMatrix_13_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_13_1 = 255'h6b792b37d68a0edcad5bdf47f1bfc9406aafeab6f0fc468237a4e28fcacbd6ae;
  assign mdsMatrix_13_2 = 255'h59ac9a2a209614991f62db483bd3908657cb8dc453f20f994954d992b9b6b3a5;
  assign mdsMatrix_13_3 = 255'h42a1ee7f6d3a42049d663211e9573b3e77f31357012971d78ea4e5a1f92fce6f;
  assign mdsMatrix_13_4 = 252'ha1c22f4712ec37852a0c375d7baba364d3896339e92a2b0b387f795312d5b31;
  assign mdsMatrix_13_5 = 255'h5bd902b72d2208f87d42df56a26d03230b2819092a57ef6c72c9e7c2f9de3217;
  assign mdsMatrix_13_6 = 253'h1dcf9a7706b9abb9214f1bf239972335d6c1e287aff618df353b3097dc6810d8;
  assign mdsMatrix_13_7 = 250'h27175b0afda75dc38e20cc8e9ef520364cbac66abc5ef762d221ebd733d7a4d;
  assign mdsMatrix_13_8 = 253'h1b00ff4ffd777d8c1abbf6fabf4365738d8be8b6cab81801bf0fe39a50bd4754;
  assign mdsMatrix_13_9 = 255'h626ad96b15dd3982031d4d2167ae3899720b157c9da6d39531359c15b041a3fd;
  assign mdsMatrix_13_10 = 255'h6a197ad26f63038b74fbef9a083571e4d84afa8170ffaf46e745208c921746b3;
  assign mdsMatrix_13_11 = 254'h349feb678f4868ab51fbe66ffcd8e6e3eee9efdfcf3e6b4a54e6e0a6f9976756;
  assign mdsMatrix_14_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_14_1 = 255'h55b1921052e9c8ea743118c7414932febe44362c3da039ff06a7dc17e3b14967;
  assign mdsMatrix_14_2 = 253'h1c30f3f31378b89066183abd44f1810edf20f4f3c81a5d4cb08e726450a52a12;
  assign mdsMatrix_14_3 = 254'h3f73fb51de0d847c4704af64bab3da3d1f93ca84a73a0660033e69a17f39eda3;
  assign mdsMatrix_14_4 = 252'h825e9ed6bae61b5310f269745dd0e0de274f6de798f94a0c16bda5104f1a35a;
  assign mdsMatrix_14_5 = 253'h1c713896047095db69cc8eaf2c2bde8521c977d7f932c8769447299c28710c8b;
  assign mdsMatrix_14_6 = 255'h56342fbbad7ece68448fc3e0f0f8c7e4b86a3b751658c1ca9ad580bd543dfe4c;
  assign mdsMatrix_14_7 = 255'h4442002f5ef57920508271e9750b87ab52d71fb71d4143994e8b84b5326249ee;
  assign mdsMatrix_14_8 = 255'h500976560cc7830e3550af4dc57e94907adde4a2c9f3b9f507c174b4b26eea7e;
  assign mdsMatrix_14_9 = 255'h49449cf10760e04fabbe8e0627a0666667f4ff3b6b9adef1f0e9d06122385237;
  assign mdsMatrix_14_10 = 255'h53c77db510957ab7b7735f477beef2af2e0e2bd28d8342ec91867535ac297af5;
  assign mdsMatrix_14_11 = 254'h32e1eddd8b9e0988d7ba042d1d80e6899b533a8411bc0782fe21f5de2e5e6b38;
  assign mdsMatrix_15_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_15_1 = 253'h199a3178a3209251b13f6b559da3e6d05fc5d182fb356dd8e7e664c212912630;
  assign mdsMatrix_15_2 = 254'h2311553bf586685820e6928b08ec5b2e5fa0275810fe900e53302e7956000b12;
  assign mdsMatrix_15_3 = 254'h28ba5262977af8b35e4fd9e4a8d762c4f3e8cb06bbf8c14dc212c44a8355ad10;
  assign mdsMatrix_15_4 = 253'h1952838952b1caea4c756a42501fa10ec630f26dce59e6a93ddc13ed146929a9;
  assign mdsMatrix_15_5 = 255'h5e7ef52923983248996c8bcbb7c2ae68db56fc4a3ed33858a6ced410aaadf2ab;
  assign mdsMatrix_15_6 = 255'h637cb6013b1ef348d2cd8327addd5adb2c06fc075d7ddf5fa955b037fc492d9c;
  assign mdsMatrix_15_7 = 253'h1bdd4ec9d45d726539e470a34e5aa34a75abd0d28ef4ac2a76c6420a94cb3f78;
  assign mdsMatrix_15_8 = 253'h17a0839248bf9a6dda2bab485ab36ba95f8fdbfae7f100b2bc3463bb57372ca3;
  assign mdsMatrix_15_9 = 255'h4e4e26013968a5236b0824c8fcea90a15329b7fad7a5f3b0119ac13b94695eda;
  assign mdsMatrix_15_10 = 255'h50e0b7a4fa12dfdd0e4391116e2749bab9b06841c1e2f9229a739072c12c0af6;
  assign mdsMatrix_15_11 = 255'h483fe63335cd025d4e3fe5fa706e764c43ac908b1574eadaf32677da489de2ce;
  assign mdsMatrix_16_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_16_1 = 255'h4fa1e46ec2c9629c747f420e68c8a02e375d636346174011b0a3df4013e5b4c8;
  assign mdsMatrix_16_2 = 254'h312e13fe6a87f7ec4ab33132a628f0f9bb32ba76fea019ddb6acb1e8145c75c5;
  assign mdsMatrix_16_3 = 255'h573591968cfdac5d5ea7c977c1a9b902bcd7d77f6e8649f09d31eddc2943c61a;
  assign mdsMatrix_16_4 = 252'hba481466b3205aa3350843a2ef38c2bb1fed57c40698b13a8137c12af7281b0;
  assign mdsMatrix_16_5 = 254'h2958476a13aa9a15a3ff4fbaae6c375bab66e1f0c8e7acab4de70f9cff5a4523;
  assign mdsMatrix_16_6 = 254'h36526efd874415309c72785e9cabd990f29f9bf7b849c556f836331f790db371;
  assign mdsMatrix_16_7 = 253'h14e788eca127f27222661c1325f6f0a76abe7c5255e4738d4b7a4c5825afaccd;
  assign mdsMatrix_16_8 = 253'h14d3d3c6394c2e2f866a6a4ec5199f5bb98979e74b074402d690e181f6ddae4d;
  assign mdsMatrix_16_9 = 247'h77eda44a4067ab26619660f6c5e7c31c7049cedc65594a3ca920e73637891b;
  assign mdsMatrix_16_10 = 255'h65907f3c4c7c312556cb1f45a947180dc1608492825ae21fc16ddf3ce8ad96bb;
  assign mdsMatrix_16_11 = 254'h308d81c4d3918cf1f073106a72ee53610505e6c636b18f797e19127b953f562e;
  assign mdsMatrix_17_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_17_1 = 251'h469a4c358545874b072db0f217a1a4e9d4e2a2b44ce6007ed830a1b84e5bfcb;
  assign mdsMatrix_17_2 = 255'h5cca0b2c9afdbe661bfd6b99d0819efaea0d99041e8e35ff2567d27e73003908;
  assign mdsMatrix_17_3 = 254'h22aa86b66e97334828e43627a114ea03e72190d239d5282a2f98c5fe1b330784;
  assign mdsMatrix_17_4 = 253'h117d9d0fea756508cce16e809d413199cd3b8725b765c9cb255a343b339798b9;
  assign mdsMatrix_17_5 = 254'h2f9e55dd0d7090e71ae4c05a8a98ec94467d5f9f4ce65e805cd5722aa2db829c;
  assign mdsMatrix_17_6 = 255'h657992b6f9fe881840bb1897feeae3dfbd9bcb3b3ce123f3ea3e43af72263438;
  assign mdsMatrix_17_7 = 255'h50f61c7a0749e9feb00da5600843852d85da8e729de0b75facf5adda984f3893;
  assign mdsMatrix_17_8 = 255'h65267370ec82496454f3bd52c3d5bf4cddc322ae8328ee952120a4af52d2a020;
  assign mdsMatrix_17_9 = 255'h4e0c97f152ac4e2be81d269ddde5c17b78ae00c61e0c2fe861fd73ee4691494f;
  assign mdsMatrix_17_10 = 254'h32d5f651b915a5e5e65352ba82e5350b2dd16055b6ed0e8b58ec072bc0a961f4;
  assign mdsMatrix_17_11 = 252'h941eb02ed99ad02fc4ddf348f5402489f5e9116551942ce722e314567caabbf;
  assign mdsMatrix_18_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_18_1 = 253'h1b392bf2cfd80b8f08761c80e311b48293883c9f97a60382131773b3efdb5fb2;
  assign mdsMatrix_18_2 = 252'he88cc2c1d560d9cdfb954af8c3f854f90fedc2a64e927839eb96647c3654411;
  assign mdsMatrix_18_3 = 254'h3d89a4dd04788448f615f8026ec0123761f60378513fc090f05793570af1b9da;
  assign mdsMatrix_18_4 = 255'h4b2d4d5ceca4d259f9e24a7332a4397babcdcc7ffd927b5c424700de5d4e24ca;
  assign mdsMatrix_18_5 = 255'h5a6e1ade0325582010ba5f17ac6fdb4c6a19dab60df2f949c8e5cddc1a6fee9e;
  assign mdsMatrix_18_6 = 252'ha519a77882a246ea31acd42f6149928236562143445a3258c642913721b401e;
  assign mdsMatrix_18_7 = 252'hfb5adbe88d65d80e3a8a3cc168e12a7467c5b8fbd265356b60faf1e56e984e1;
  assign mdsMatrix_18_8 = 255'h4c3435316760ed635aaba8cb76db9b22ef4ad135a050d60bb6f073f493e3e53b;
  assign mdsMatrix_18_9 = 255'h5ffa83810b5ea238bdf860e4f6bd77182822760045f81e462df7b35dab4b63f5;
  assign mdsMatrix_18_10 = 255'h5910281b6f75f951a90eafe4dcf7f6f45f28366521df0dff84913fd2b797046c;
  assign mdsMatrix_18_11 = 255'h694373266c05a225c23d2d749e38ee9c914d1b5dbb2e197808ac3f056ddf4eab;
  assign mdsMatrix_19_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_19_1 = 255'h531d2a39fa79f939d4cd70793107ea5d346bc1d200ccf532a25f9f3a33cb6b7e;
  assign mdsMatrix_19_2 = 255'h49fa548cacd2ec82aea7ebf1d0254dba077d45e3093227e955e1dbcedb6de606;
  assign mdsMatrix_19_3 = 255'h5a89b30789a923c20148c96f531dcefd96efe121a211fe8e6586b871a364185d;
  assign mdsMatrix_19_4 = 254'h3ecd161d8096c0f1930e541ca70aa5d2e1c18b7ca2aeeaffcf98c02e1bacac60;
  assign mdsMatrix_19_5 = 252'he96ecbb128d47061bcc1825b3d0f5e85ad6484cb2671a6e88bb0db1c5b6840d;
  assign mdsMatrix_19_6 = 254'h38d20dbda2b7ef8cc8044687b51f0558a2dedb8ac82d97a01acf43a48248b1ea;
  assign mdsMatrix_19_7 = 255'h465fa699babec84cfde035e90c2e512c705af5acc6f4823f36887ca5ee48a53d;
  assign mdsMatrix_19_8 = 253'h184f320bea3c141058275b0bc91e00e49a2c3ed5e3ba38ad5d92f862eb2d0408;
  assign mdsMatrix_19_9 = 254'h2a06048b9ef62cabd11f6f113de8b58ea0ce2baa42bd7e9f4528efe3b8c9112b;
  assign mdsMatrix_19_10 = 253'h18e6b3df871f150ec4910ffb4da47a3dd1c0bdf3464998e4e8178d5844787825;
  assign mdsMatrix_19_11 = 255'h735a069ba4eaf2fbecf3e9414b625705985904146965ff71d2a8a1de3f0e0823;
  assign mdsMatrix_20_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_20_1 = 255'h69327c13ee54509a355d5a92aad6566ff52b4272db544dee0f63adab6c051b2b;
  assign mdsMatrix_20_2 = 253'h14ebcda72f4d7e2a863b30b8aa58b8132e00590c7c107103b412c317b4a9f4e0;
  assign mdsMatrix_20_3 = 254'h2b1e6fac4b4a8d9dec9c14d4515b9e1aae95513e3f021184696a6258a5716441;
  assign mdsMatrix_20_4 = 253'h169d54c34b9ed10117c2fe8c260cf04217273498110ced3eaf88f1c30b629a8f;
  assign mdsMatrix_20_5 = 254'h3d00a07f349e95934f44d71cdc0086a277bca342cf2a38e9ad1757150d490191;
  assign mdsMatrix_20_6 = 255'h45a57dd3b77a69c6fb9d69962de76d9ee3ca2d8ab141203b5b0ab29b14c62491;
  assign mdsMatrix_20_7 = 253'h1984a3e49f2466b69bc6117c169bf408f1e58f259e4e2685c1fb1cc2e0e6ea8d;
  assign mdsMatrix_20_8 = 255'h565c811ab57896ecae2b6049ccdb113fa7b9faf52374633febb5e7caca766800;
  assign mdsMatrix_20_9 = 252'h81079d2b950216161100c139dad2c796d2636fa54577fcaddd9f024e1fb31e7;
  assign mdsMatrix_20_10 = 254'h23d2a4f3d52eb524e9f98e67fb897f4233b6b7c7328ea0b19ac4e722109166f4;
  assign mdsMatrix_20_11 = 253'h1a48fcc0921ee76b4231fe75b239a3c846c48f76d86c8b94e29473f985d14d2a;
  assign mdsMatrix_21_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_21_1 = 255'h5ffd9ed4fe6d1c89c3cfd88641b9a6d65b198520cfff9d5209d50e8144ef75dd;
  assign mdsMatrix_21_2 = 255'h49581a39baeb2f971b4038ff7842ec267b97b05a063008954fe544176c27e205;
  assign mdsMatrix_21_3 = 255'h569193badee1d4dc2639e28bb48cac7bc822db9da7f2810d43386136fb364bc4;
  assign mdsMatrix_21_4 = 249'h154353d9e356e3755e20e3854525059d53867bd124e5c531d3c3f6e10b4a2c4;
  assign mdsMatrix_21_5 = 255'h4a7468d8c153b2a91692d008bf060d6437f9a8ff897881a9e0ef3a212cfe671d;
  assign mdsMatrix_21_6 = 252'he36bfcd6aa4f8044a0d39b3fbedf0b56b6ff9c2769d881c4c3012c219124511;
  assign mdsMatrix_21_7 = 255'h467c742c6d5775917a4e0ec3d1eb9ca47ffbf4b06b09279594f44afe5b06a733;
  assign mdsMatrix_21_8 = 253'h1085b21dc1ba1a19f5e5571a858622f34baa0893341fb0ce70e6269347c9b4ad;
  assign mdsMatrix_21_9 = 255'h584f3983e1684b9cdeadc85e51367c9207e95229a56d5a358733ccb709188d05;
  assign mdsMatrix_21_10 = 255'h45c3f6f6b3fbc8cce98a3098dc21b808cbee4b5024b0939eeecd564cc1197d6a;
  assign mdsMatrix_21_11 = 254'h3c62554a8e1bc8f352a760f488a011ee5fe3f60a8140a1b08d3f6c99148e84d8;
  assign mdsMatrix_22_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_22_1 = 255'h406c385463c54985133c96eac37247c908119ff16a84c0e04f51ffaae966e684;
  assign mdsMatrix_22_2 = 255'h6a6f0287e6fdb3953bfaaf653a8867a08ead9c42e09c878a593d827021484621;
  assign mdsMatrix_22_3 = 255'h5f34c01f2b035db4f87890037d97b0fca5ab23f912b021f5761c3b6967f9d423;
  assign mdsMatrix_22_4 = 252'hdf335bc9326385e1e1a62ea3bd5315b7c9ab13f3aaf37a4a45601fc13959ac0;
  assign mdsMatrix_22_5 = 253'h129cfdb7e4af2a1ecb48ec06e46cb1e9bccddc59204d5a687510261f47a53bea;
  assign mdsMatrix_22_6 = 254'h26aa973699e1c36a22577c69c67a4b93703ca30630a5c43b8f95a1b66f04b4b8;
  assign mdsMatrix_22_7 = 254'h28f320fad070b6b3e4b483c5f0d2310df9739d7359b5d467abd4cf2514da9121;
  assign mdsMatrix_22_8 = 255'h483437e7a3a10eeaf55dc709f05ab886833b0cdecdb42faab798fc078d63cc4c;
  assign mdsMatrix_22_9 = 254'h2c1ce5458b776fd46523648212a63bcace53ddf82193fcf65c771e920a29e060;
  assign mdsMatrix_22_10 = 255'h42ee234d15959540da48d8cbc15b3e935917309d7ade9c3028ee2923b405a297;
  assign mdsMatrix_22_11 = 255'h4f021b3146e2ff6db986d878a07c01bd6619917b5335cda038b005e010006d8d;
  assign mdsMatrix_23_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_23_1 = 251'h7763d29763a1238e0894967f76515c37afe0da6ba940c8028b0bef061e22494;
  assign mdsMatrix_23_2 = 252'hb907b67f66ea6be26df06bf059c95a39988dd509990bfc5d51c95c34de3cb60;
  assign mdsMatrix_23_3 = 253'h17bc5e5f13fc3446d3d66f413681b9132ea4f4e8c0230b3d8ec64719ec055b61;
  assign mdsMatrix_23_4 = 253'h11eeb98db9e00eb7d1b2f3b5114d53478750dd4783754f052c6d9de8732f8b65;
  assign mdsMatrix_23_5 = 253'h19addd67fec355b2880cf2c4bb5ad89c7634a5ec6c6abedf279d191e7cccb5dd;
  assign mdsMatrix_23_6 = 254'h2dd902b7142e54c217cea3001610d8a71e962403849c454864f19c41b3161aeb;
  assign mdsMatrix_23_7 = 254'h2a3b32c4b36d3e4775f193577ff86ca2916ff0873e40a5d7f9f557ef6f089dde;
  assign mdsMatrix_23_8 = 255'h48fbea862f330ba77e5024cc13b6e4a15211a726cd24a48325d5f61cbbdde0ae;
  assign mdsMatrix_23_9 = 255'h6aa4b6a67a89732ea39cf3520f293762b021d575708b6f1c31d48e2b4ce078ae;
  assign mdsMatrix_23_10 = 250'h29c251880f45b7025824d49bfc6594a74dc53e2384354b0c9ba974cbfa1d406;
  assign mdsMatrix_23_11 = 254'h37b657bc4221a606a9234981e12f4208c4a666f250739537a4188bdd488522f5;
  assign mdsMatrix_24_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_24_1 = 254'h3c1098b26990fc5e89e16581e63f80e9c1c471e379d9a635f2684da5eb86c800;
  assign mdsMatrix_24_2 = 255'h47f2143f98ffb7d503ab21d84b482cc28bad359df4ecb071b7a2650823ec2d1d;
  assign mdsMatrix_24_3 = 254'h3c43dbd9befb1111f4c894205ad14625b78f0c2045987e9c50216cd3f391c4ea;
  assign mdsMatrix_24_4 = 252'hb3bed16b04ce040f08b4c1ce9dd28cb12be9318af456f0fb050ab3cf5258641;
  assign mdsMatrix_24_5 = 255'h42f69075f64eb70779608f3d1157d03e659444001fa3d01a66aa8b292fbd1029;
  assign mdsMatrix_24_6 = 254'h348a77080c56dee1dee930673a92510e38c1a317e78ff940787d8cb56100a174;
  assign mdsMatrix_24_7 = 254'h25ca0831f008674cbc24c6ee1ca6fc0ae27957e6d70eb3a1a15b017cf64f4e6a;
  assign mdsMatrix_24_8 = 254'h36a37be4e4869bbe7fff897d427863e66682e1d78c1bcda777555202e1e1faa7;
  assign mdsMatrix_24_9 = 254'h256f7e1fa33843eddc6422abebb3c37da362e793ea193b6b2e404fb5d6eb3ec6;
  assign mdsMatrix_24_10 = 252'hd511c9928a1b772a3a176f0d703a9ea8b4892df0a7b73748ebe1089c05175a6;
  assign mdsMatrix_24_11 = 254'h2e74ccafb35c2c5090ec072e303a310702411bd4726a6e5eb58b0eff3737c826;
  assign mdsMatrix_25_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_25_1 = 255'h4ac465824227afa3c57542e9f8a0e4265ebed3ce155590bccfcb709bbef78d92;
  assign mdsMatrix_25_2 = 253'h122c47d1e327a40f09cc0ee2b89b3d200c460423e9843564dd7f18dbca652166;
  assign mdsMatrix_25_3 = 251'h5744c936dc179d845c05b70fa9acb5882fd11babb611d3fb2133fd6b83ffd28;
  assign mdsMatrix_25_4 = 254'h289e08b17ba5a133c43a53dfa8b29fa19f044df82ce7816e36c40d566ef48eb5;
  assign mdsMatrix_25_5 = 253'h109e679f0032fa9e8db4c88d2463c66ac5fb1967463ab414071366b904c122f1;
  assign mdsMatrix_25_6 = 254'h380e2d02c016438e0072a64e033ce14a495ffa8851a5e5d64c78968a41bc1c59;
  assign mdsMatrix_25_7 = 254'h2976d5373eba54dcae919e191bc439b6d262a6d9ebdbdb8d6bc05574d553812d;
  assign mdsMatrix_25_8 = 253'h1bd89a08c76bc9f656371e0cdf45493be3332a9cdf47415b419f1d27983953d1;
  assign mdsMatrix_25_9 = 254'h303234db32a95d2c815302d7d3b9cd6394794584f51cd00df176ba01267d90de;
  assign mdsMatrix_25_10 = 255'h55ca8d9a14849c36d4a62939fef8095cc77a3c278f3ab4bd582e2c1360548194;
  assign mdsMatrix_25_11 = 255'h4889cd07fe76c275d1025625faf90faff0c00c399a27d7a287a9bdb3dc6fa28b;
  assign mdsMatrix_26_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_26_1 = 254'h3793fb86de75f82647866c61a9c3af113db61be4591d73c3561728b9631e09db;
  assign mdsMatrix_26_2 = 251'h52cb631538544c3649aae29d7e10d5620b458e088eecd59e37e6de90a57ec82;
  assign mdsMatrix_26_3 = 251'h60c7ccb596de9b44542e373a6f3d9e633e95e177742fddc8533d044c8858b8a;
  assign mdsMatrix_26_4 = 255'h59633d7eeaeb1a0620d7ddeb6024ab7cc98a180d4b45fae6644a3295d5f9eaee;
  assign mdsMatrix_26_5 = 254'h3187ca8aab4adc634e472f35ee1aa08bb77ad8fde8708aa778137a4dbf5176f9;
  assign mdsMatrix_26_6 = 255'h4caa27f8df02127b173a7ce4f05c8e94217e9d988b3da6bdb8ac5f5299360736;
  assign mdsMatrix_26_7 = 253'h17929124621b43c3e51cce8536a882c710e5ecf664317cc8f042fbf6d5c46d89;
  assign mdsMatrix_26_8 = 255'h5eb91977f5851528484a3a552dbc603935e38b2bcca607fcec668980fbe1e4b3;
  assign mdsMatrix_26_9 = 252'h989679917ccf0d7305923c2c362b2b85d4aaa111a0fc0501d1e4c7d7c783aeb;
  assign mdsMatrix_26_10 = 254'h213622df17ade4abfcfc785b71f30621bc03b09eec4b5beab08390524b15a597;
  assign mdsMatrix_26_11 = 254'h3fc23e71a05a531c177d889f41085b2cfe37a22b7ee610bfdc61716d49b6ebb2;
  assign mdsMatrix_27_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_27_1 = 255'h68bd4a7c62a25b2a5e9def071fed40e5a5f3cfe0205b55fd03b258507dca77a1;
  assign mdsMatrix_27_2 = 254'h29960eece812146c4489ec6315de4e2b7b9db11a51cacb926819ae9a337498d2;
  assign mdsMatrix_27_3 = 254'h38fdc599d85f0400eedde3c8e0a55bec6b147fe9407a67d790000ee9c3c9be55;
  assign mdsMatrix_27_4 = 255'h64472e3f075c2319a230af10c826aa742cdb116f2b962ed23f13513ad40ce1c0;
  assign mdsMatrix_27_5 = 254'h3f3ac0ab959748d3afddb4386796aedb6d5625b7fe417b8646375de9d551edf2;
  assign mdsMatrix_27_6 = 254'h33715842cc55a41ad2bab044c8b9fa04fc3ee23264313f64413cb14459c63fc4;
  assign mdsMatrix_27_7 = 255'h52eb2616ce640592c933149ccebf5ff6bd50a4b86b4aa82134782e0dcafaa4a9;
  assign mdsMatrix_27_8 = 255'h50fa7cb1d047a87b8fb2b5a88398fc55bf8ef59c4a17b1d989e680c3a2443097;
  assign mdsMatrix_27_9 = 253'h1d0bbf3ceea28de6afad2a52ad1bfbd97ce8ccf74684afbe8cd0d2e80570edf3;
  assign mdsMatrix_27_10 = 254'h3b4f66280d49b308c85425fec134f989ae106bed9356a50842d6bff0ad34a6de;
  assign mdsMatrix_27_11 = 253'h1fbe4c8a3f77a4025e79b7eeac64e82be3533de46945cac860cb8891564999cc;
  assign mdsMatrix_28_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_28_1 = 252'hf83c718ddbcfc638e49715fcb9df2360052c9175ed16b1739b92473a566a5f5;
  assign mdsMatrix_28_2 = 254'h33a430287090fcd9170ffea2eccdc4f65beff4b77c26f3a6bf2f493b42d91397;
  assign mdsMatrix_28_3 = 255'h6bff8f4505fd15722e7aed2c4fcae4f101a7901478341bee15cd29c41d43509d;
  assign mdsMatrix_28_4 = 255'h40fed8c3d8987f149d4dd6efa445e2ca5e2972402be325c1f224923a8edeb5f9;
  assign mdsMatrix_28_5 = 251'h5695855b7cf9940f734a1c5ea924aea7bcab5ba3f48abbfbc4669b2fae92905;
  assign mdsMatrix_28_6 = 254'h21daad558b085c2a46f201f88e7a9622f6f26f7fbeb59790705439a7201281fe;
  assign mdsMatrix_28_7 = 255'h47f902e4b7bbb2bafd4de2caaed8c9bfa1614bc30b5fd5bb80d3cca17d77a06a;
  assign mdsMatrix_28_8 = 255'h668b12d059310884f96d40d9193bf7dd2d0683f23e17a98e861525fa021d7da5;
  assign mdsMatrix_28_9 = 255'h5e021cbc30fe9129175f467f802810322caf71afb7d4563d5eb37e92f54f03e9;
  assign mdsMatrix_28_10 = 254'h3aec6ad41c6a63b9f5bc1117ba19e1a0f1f0fec90d0ed9113b04a2c1188ad896;
  assign mdsMatrix_28_11 = 254'h259b079b481fa135b77ad461df38cbfc9aa8348f8a50b866d1adacc940ec38e0;
  assign mdsMatrix_29_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_29_1 = 255'h72565d5806f9184b76220ec1da98f4cdc3215a6df68786b82cfb9f3bf0b6f28f;
  assign mdsMatrix_29_2 = 254'h22b6614c59b3994f43ee4e3446b48aa69a6c12e22b6b1a5ba6225caf13fdbd6e;
  assign mdsMatrix_29_3 = 255'h4631d9c23c2d31908e1813465f241183738e6d62e2baba5654e35b13265bb702;
  assign mdsMatrix_29_4 = 255'h6d4e06cbbde6444ce5da5952bea53fdb5119d6f254c7062436829e752ef06902;
  assign mdsMatrix_29_5 = 254'h39a23cfd6344cac87c2f391da86c63b5d4788b5c3ae0821e0305565e3a1601d3;
  assign mdsMatrix_29_6 = 255'h66617547b0e8a66a1fd48112b3220c5a3ec668b4305924596e5ed75f2d4ffcc0;
  assign mdsMatrix_29_7 = 255'h44e66243e7316409bff55b2621a28609213ca68274a0366992f486d7d43fa6f1;
  assign mdsMatrix_29_8 = 252'hf5fe97f7e729ff4f2982dcae31d6612571b49b26323cef74563451fd1d28c18;
  assign mdsMatrix_29_9 = 254'h340142b8b203faf625e319ca0f6c759aa3edc782280bf94288f87c26fc8b7a40;
  assign mdsMatrix_29_10 = 253'h15aee466606a483bce3f1e8939bebbccc89fd2ed2b93ad41fdecc1cae56aca82;
  assign mdsMatrix_29_11 = 254'h39b4544faf6775ec2a7cc9b36001296de52d014d5ce4120971b96aa506e6c579;
  assign mdsMatrix_30_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_30_1 = 254'h2acc635f48293a4b20fde809978503d25af46d3e6c471e474d62c00de2de8c77;
  assign mdsMatrix_30_2 = 254'h326f1ab03a73402ae2a4dc8587ac46e999dd93b16b72f203deb30a985c3e94ef;
  assign mdsMatrix_30_3 = 250'h37105091adb5640d30ac6d1d74fac4df1f604a7a25ac2b31ebea5217c22669a;
  assign mdsMatrix_30_4 = 254'h2b71a69ea6acd614b64d2f39c7f7d67e1fee6c93330bd179bd87511b748855fd;
  assign mdsMatrix_30_5 = 255'h6d9fda4b6b65ea326395d56595564f96deabc6e0a5de68c79af20bb80c8d47d7;
  assign mdsMatrix_30_6 = 255'h50f197f9f021f15a1d9d9a893f55f3e8c96587ff68f3e7791ca07141ab6da1ef;
  assign mdsMatrix_30_7 = 255'h4ce0c80cb05ae39f74ad0aab1c83173704f3eb722fffcb87a4891c2bb95a182e;
  assign mdsMatrix_30_8 = 254'h3c8cfa1c32f28c2ce8a487d077d303322db47111275b94526ae85d0a2083bff1;
  assign mdsMatrix_30_9 = 255'h4cd5df61f09c86212297758eb8e7e3452ab57a07bf27a9440cc93cb02cd3c697;
  assign mdsMatrix_30_10 = 255'h732ceee618e067d1ef76112ebfac5d8aa56bad5baf1cb24ca962153a5db7bea6;
  assign mdsMatrix_30_11 = 253'h108681cc424a4e7d59bbda0a8199004e4db811b3e91d45dac8b6723d245fdee3;
  assign mdsMatrix_31_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_31_1 = 253'h18ea9199876ad6edca425c6b320cb4b6d159ade165863c15d05f1f41c579064b;
  assign mdsMatrix_31_2 = 255'h6701eb9325a8f44059d6d093291c5ec1aea6fe987623acc49c0996f30acd393f;
  assign mdsMatrix_31_3 = 254'h337bd609fd6551583f1dc28be28cdd438a7ac6f32801db3f372ac1447eb2c7e5;
  assign mdsMatrix_31_4 = 253'h163ded56a8aa783937ac7e3ab98fcda5ac08921cc9bfe8ee7b314871ac1591bd;
  assign mdsMatrix_31_5 = 255'h5f9c0773b973cebfe16183910ec62a28f2893b87647207b256f4da1d1b74ba9e;
  assign mdsMatrix_31_6 = 253'h1d31f34393f4f346146ca380ce843e70ae71c22dff1add6c054f3f48e2d0f5d2;
  assign mdsMatrix_31_7 = 255'h6c8eb7cd0e8c6cfe34675926c7835a219a870bc51bd686bb97d16007f2665900;
  assign mdsMatrix_31_8 = 253'h10bc3d55b87587b511ce4fdd70dbbe32b2dd7c9d6abb090fd8e2c02747b89f5c;
  assign mdsMatrix_31_9 = 254'h2568edad66128909f42aa8009cb50f3db68c6444524251bb6d76fffc3d827f69;
  assign mdsMatrix_31_10 = 255'h66d7b412102e4121096aaa3d72fd4692a48660e917776a340ad5dfdab6e99d57;
  assign mdsMatrix_31_11 = 255'h5916cdec8cc697c6cebcbf836b4eedc3bd96ee60e347064d7eb7a4f59e8de3c5;
  assign mdsMatrix_32_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_32_1 = 255'h72f1278bc7e49af310205876eacbdf32b0ef97e1fed1d32412e13558678b77cf;
  assign mdsMatrix_32_2 = 255'h6e6647f8dccde9dd8d35aa77202bf966faeae511cc36c66ecf418048f11d9240;
  assign mdsMatrix_32_3 = 255'h5b95a5661fa7e769f0bf383d888eaccb99e13fceba3527c96379521f1547ed5f;
  assign mdsMatrix_32_4 = 255'h71da61f99a73fb62a3cc09b273b4a6f7e963c70c4dfa4e390d8c8a6d88ea460b;
  assign mdsMatrix_32_5 = 252'hf3c0df2f265adc840ec856f7715ed12c754ae2c2272b7d1477480f675687847;
  assign mdsMatrix_32_6 = 252'h91e5aac1a09b8ef5da24844bffed1ef2ff8c98d489df71fcb07bb8d1188ecb6;
  assign mdsMatrix_32_7 = 254'h32e56332427a6e69086ca5be3457d500c6ed8fda1c7823f391be0031c0e15e20;
  assign mdsMatrix_32_8 = 255'h5ff64487227be1360881f631795d00730b651ee985068bdf7aff93e5e33ee4d6;
  assign mdsMatrix_32_9 = 255'h69bbf6e9ece39df4e02d181be1b046072776bf9e5b9e49581757508f1f0bee6d;
  assign mdsMatrix_32_10 = 250'h34149381f7e94f0e5bbff63e320d978ab2a7634891129dfff5edbef9ace357f;
  assign mdsMatrix_32_11 = 253'h10b69a29058f53e989ab27cb794924dc51ecfbf04a9bc2dbbe72428291e1570d;
  assign mdsMatrix_33_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_33_1 = 255'h6dcf5691bb1619c78bbbafaecd92597ba6412c2111eedabbe2a2bfb09b80887a;
  assign mdsMatrix_33_2 = 255'h5961285ecf2fb49188cb9b46e64784a78422a4c2b74f86e2948cc0cac7131646;
  assign mdsMatrix_33_3 = 254'h22a856e102db10f50dfef155d77f439e0b918baaeb473c86881cd4257bc36c93;
  assign mdsMatrix_33_4 = 253'h12e0ade4fe058aa7a943eaa6d055ca820c03b9d0a95217b5d8934a7e5a544ac3;
  assign mdsMatrix_33_5 = 255'h64af92daca652ebc682104cfd4a65547adb8ae998ce64671f3864a1ba486f69f;
  assign mdsMatrix_33_6 = 252'hdedbbc3556c64c46605bb08a628df93c520e57c98b743e923bf94be1ac3974b;
  assign mdsMatrix_33_7 = 253'h150fdcd22ec031baf30108db5e2cc1aabc9a18760afe752b1f6a6831b1b78b00;
  assign mdsMatrix_33_8 = 254'h39cb2882d32c761b490e61e9d4e11c86fe029dda58f42fa45fe764004b2bc8d6;
  assign mdsMatrix_33_9 = 252'h8cdaf436f2355556e34022b4205b45306544289ef8e2e739a50feb93d45f095;
  assign mdsMatrix_33_10 = 251'h501c8316e7a4f09b784537eaf99f75f1935abc7862bd0409442253ad46dbeaa;
  assign mdsMatrix_33_11 = 252'ha1c8c323ad47611acfedc69952c011167bfccc9ea717eaa3dd2405052878cf2;
  assign mdsMatrix_34_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_34_1 = 254'h281f62947f2da3a40183e73ad3bf7efbbedd597302c92564515541fcbee38b5e;
  assign mdsMatrix_34_2 = 255'h46f64dfa79531097bfea758cd1adce7e3f3c3839d268a1723286274ca082fc41;
  assign mdsMatrix_34_3 = 253'h13e162a1678b299dd182288b757b55f68ab769e01fae935ddf6a93b6f8ee73d6;
  assign mdsMatrix_34_4 = 251'h7e9dffaf1b9ca8c7625b299619163192ce4d2b876306b07f9d4efd84d8bf60a;
  assign mdsMatrix_34_5 = 255'h5c3fb47686c84ec67caee4fa1d2f67b1e4c8d14a73cdfefb3c49d3da1fb12f1b;
  assign mdsMatrix_34_6 = 255'h56bafabc3f4363e0ca6683d40f06a061cafea6df1dc7519f675599dbfbfeab1a;
  assign mdsMatrix_34_7 = 255'h4eaa0cbb2bdbcda42c81763e1138bca132e3b03af76952b953bf9c78fc59c513;
  assign mdsMatrix_34_8 = 255'h4bae10d67d8ecfce04704405077f39a6bd3daf8776cfcda191f149ccbfe46704;
  assign mdsMatrix_34_9 = 254'h2fc7a9cae3eb7295a3a7fc3f5e319915790e1dd1610f82e1127330d807ef6cef;
  assign mdsMatrix_34_10 = 253'h1d9a46adf8454445d4728b72ccbd9531eaa133cee645ca4477ffb1a2e157fbb6;
  assign mdsMatrix_34_11 = 255'h6d3c465713e5ea15cd10425ce79ee3da7395cc7fb3e835902f01b562a1d246a1;
  assign mdsMatrix_35_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_35_1 = 254'h3d664f8b584591db73198e2dd4e5e81d3b1f61a2a67b02d1d09443c6ee6ecdf2;
  assign mdsMatrix_35_2 = 255'h5e0f417cebad8f8a43d46caa20d33113213150680fd3b7345ea4daa18292aa8c;
  assign mdsMatrix_35_3 = 255'h6e2bae1468016feef59238d07e4e19caaf4fa629d8eef1fd46d1fc7cb55963e0;
  assign mdsMatrix_35_4 = 255'h61078da5839d88533f950c78fd4f12d1f4862723e62c9870e4f5b76dba92f02c;
  assign mdsMatrix_35_5 = 253'h12fbfc6a07d437ca504fb6d518164b3abf8cae5be5fab256f9ec0d8bafe7a9d5;
  assign mdsMatrix_35_6 = 254'h3e6c460421f0f641ebe273ce90a979d5a6e6b9cc5d35e302816372b90e8e74de;
  assign mdsMatrix_35_7 = 254'h2b1b1f7e9cde4d2b8670e76876d1d6e981d19c568e7c7757f3b27bd9733e2dfb;
  assign mdsMatrix_35_8 = 255'h63fa6b8e824a148e6375ea9899e86804ca9c39ad61f048c7f49667fc76f13702;
  assign mdsMatrix_35_9 = 253'h18e39c371056fa345a8601d8a75ab7d7cbaea9403cfec402aab940d16a2a6b38;
  assign mdsMatrix_35_10 = 255'h600eef4f6f8164f7cf3333ee1ccbec655ecab62fc7f0c72015059e9d5083bd5d;
  assign mdsMatrix_35_11 = 255'h550fe6d38ba9b7005151950e82b3f60e8856bd4f66271c9dae34a82ea8911e53;
  assign mdsMatrix_36_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_36_1 = 255'h699558ae99162096a65f8400089781ed054a63739177c641102c57faa82b18a1;
  assign mdsMatrix_36_2 = 253'h1d42c3ad0cbf0d7e27803a8d111028f792864f78006526ee6b3c05f74a11d42c;
  assign mdsMatrix_36_3 = 249'h16744ba8ec7189364b2c8930ebec036f92ea0fba1610ec95dfd07d211258e25;
  assign mdsMatrix_36_4 = 252'h9c335c644f977263f2a26899c15880319c2da63212b9fa8c8bfd7052810ac1f;
  assign mdsMatrix_36_5 = 255'h6097ce819240c8acd21e9268784af92bd1c2a66b022ff8b9e8b7b50f319bc084;
  assign mdsMatrix_36_6 = 253'h1ff7b01d73fa76ba51db99dac8be04ee231f71a68d7814a5cc9ad1457d677bdb;
  assign mdsMatrix_36_7 = 254'h32f1ee9ddcaff76e3767c9e2462c1dd969a99deaf4869db9f9819880dee782bb;
  assign mdsMatrix_36_8 = 254'h3310432b7d739d37603fa2e2bb822b37e2a698a8b781967ec355ada4b2a59cb0;
  assign mdsMatrix_36_9 = 254'h28ace45a60c1a5c259ef474f920f20001f0ecd10a818468e5c7c3b4749a42cc5;
  assign mdsMatrix_36_10 = 254'h2df464a48901e3d65fec6167a82d9b4f5eec4b8d1beafffa963492eff5a6dcf6;
  assign mdsMatrix_36_11 = 254'h2ffe7f5a1a913651ddb666272acf7555f82c60b3b6772f2d74f570d6c05b4685;
  assign mdsMatrix_37_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_37_1 = 252'hb26b95ba465ccacb8e6953bc4c04617ceca07c39fa12feca7d130c90a33d086;
  assign mdsMatrix_37_2 = 255'h47df322ff238f1798e5f4df1252f6973d7f0961cc562a39efd018241d79a9be2;
  assign mdsMatrix_37_3 = 255'h65944a0f9e38384a8d693e9606c9fe251d6aa5cff52082f40412d6c596691032;
  assign mdsMatrix_37_4 = 252'h94b73ce679592ec91517776b35fef6deac7e4dab1ef4bd2e3586ba32e010db9;
  assign mdsMatrix_37_5 = 254'h24aa3066c26c022b6789394e3d494f149b1c2225f49b538cc87c67f7932a8fc9;
  assign mdsMatrix_37_6 = 255'h442e25ca2b98a24e6edb093a7e28a7ab1218d1f456fdcd17af686ecdb14c8219;
  assign mdsMatrix_37_7 = 255'h68d7305180fc0ab4135b79ed77ab0b496665390a3c19b9bdf07057358972376d;
  assign mdsMatrix_37_8 = 251'h416022c39cc9f04577f5239e23d365f5d89314b966d8633ad9b7280c484f25d;
  assign mdsMatrix_37_9 = 255'h4faf22b3b2eda8f055c4f2d4f52ceb90e7494142c2e38000706b8d55aa98ff6c;
  assign mdsMatrix_37_10 = 255'h50fc8cf24c32fb627693eb4bdf7ece6c360ea4022cac967b7ed6b73210b92688;
  assign mdsMatrix_37_11 = 254'h338c3b33348bacfd9dc66db054f4792b0c693bd7bf650c407a316da763a931f4;
  assign mdsMatrix_38_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_38_1 = 254'h3eee7ceff58819a1a652a7f26c9fb47b004e87c6d21be6722bf515fbce1f549e;
  assign mdsMatrix_38_2 = 255'h495b26b26aa7bfe1f4a1378b135a7f14c58751edb1f9056c4ab6ac34805f4523;
  assign mdsMatrix_38_3 = 254'h3c3facfe1570e84d72288947f1f2db353954cf97d518cb143af03a9ab5112dc0;
  assign mdsMatrix_38_4 = 254'h25a7aaa04a875f528a3aae78df5c234c6226b6281688b377a528c3fc7f4f64db;
  assign mdsMatrix_38_5 = 255'h62e7db1984b4afbeb17c1b36f03718b493866401f423b0ed60b36c006ce59345;
  assign mdsMatrix_38_6 = 252'h9546d516d02651b9b766bfe1bcec37e05dfec5905dec84b3bfce29b65ec4903;
  assign mdsMatrix_38_7 = 254'h22a78a397404f592ba5921cfcdba4b1997586980bc9d054c98caaa7b29258f6e;
  assign mdsMatrix_38_8 = 251'h6f5ca89293e408a1e886c2b3e8451babd133026938e8ff2b182b949b0e6c05a;
  assign mdsMatrix_38_9 = 255'h5501e00551617520135b771a6b3e8929f28ead8a62957cd555a2590acc8a7ff3;
  assign mdsMatrix_38_10 = 255'h66f260b0c42df3978c90be7e056718eeab6495749bb21e76ce837152ba0e184f;
  assign mdsMatrix_38_11 = 255'h7340b475fd1ea09b08839ec216d18787b866fb1df9603789f23742863eed4036;
  assign mdsMatrix_39_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_39_1 = 255'h4ae782de2c3d7f431f1df5e0f95bf2a372a05f4d63852a06f2e70e1fd85e676f;
  assign mdsMatrix_39_2 = 252'hd21c6514d14a3401554c7bd041ba6733cb6241cd9a76ab9398c831845ed8944;
  assign mdsMatrix_39_3 = 250'h37910621b1b0e06276a34a3d4845f12aa9da4dd9c6bc4ef0b6509ad4482b7a7;
  assign mdsMatrix_39_4 = 253'h1a65b567de92bdb40a04cea84320809f6677105d884728acd87bcc5a5b5c84ce;
  assign mdsMatrix_39_5 = 253'h19429d4649329c9a1aa6baea8001dfed0b1f837e35d09d8e500086fd5af2cca8;
  assign mdsMatrix_39_6 = 255'h726068b843c0044e4280886100a245cdae659de2019f765df762c37fd62924a4;
  assign mdsMatrix_39_7 = 254'h2dec9ab28804210a09220608f4c44bcbadebc1291ed6d4fa899e479a999271c9;
  assign mdsMatrix_39_8 = 255'h5a811f58377b553d749b389fa3079d3045999647e2f02ad46b7a409beef961dd;
  assign mdsMatrix_39_9 = 255'h46cf8f4663d997c4708df61afb62d8298d977e047c2e4097252236be2a181884;
  assign mdsMatrix_39_10 = 254'h3d14d717c5d6fecea7e576cb57f76fd39a4ab25af2f9ae4f5909013cb4a0fb34;
  assign mdsMatrix_39_11 = 255'h6acdee8e43349a392c2dc80fd4a2a58736bddad4a284dff4d64974cdde20ba75;
  assign mdsMatrix_40_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_40_1 = 255'h596a2e28089eb4b0bb699e63714a7cbd13dd33f8a1f2808a75d0d081a4b1fa98;
  assign mdsMatrix_40_2 = 254'h3d950e5e483d162f563e95619ada29648ac924b3848cf1710a3e4e1549e5535b;
  assign mdsMatrix_40_3 = 255'h6cecad8af46a9ae7c4fd6b2b6b3483e8c8b94ab5d4314a6e3d6b4497ad51cf64;
  assign mdsMatrix_40_4 = 253'h108725ac41951acd5f796f78a550917cc5d78f999bb166cd16d8045d3017b8dd;
  assign mdsMatrix_40_5 = 255'h529c31770a594294595cc91aa7ab7066d441851e34fc4906e9ce75efe8b18cd1;
  assign mdsMatrix_40_6 = 252'hecd4e5e701a43b4482fba24aad7749e154f1a932515f9163e5e2a58ba052de4;
  assign mdsMatrix_40_7 = 255'h5cb43247563c5b2055e493a50ebd1e6d18210517b7f2be51eb5c7ea1ebbe1bfa;
  assign mdsMatrix_40_8 = 255'h6cb7cb7911c47df5e8021136d592fa6b55f61e2786fe793855c1b1bce879e870;
  assign mdsMatrix_40_9 = 254'h3a4c8bc5b366c15039cb506a29abcd880c6d18b03e2ce4dee928b41cf22d7d14;
  assign mdsMatrix_40_10 = 253'h15da39c9db23d979fb60d29a24a0fc8c2e2e3b7ea2af0b111cf21de2e78723c7;
  assign mdsMatrix_40_11 = 251'h5f243e47d5111c185d11585b1b0b9577aa8aa448e460fde1d70217bdb2a6ef9;
  assign mdsMatrix_41_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_41_1 = 255'h456802388e41176db5cfaab1e9c85e61ec688bf2a9807ccf031ca68f4adf1d16;
  assign mdsMatrix_41_2 = 252'hea567d13f45aaf978adccac93e011a3a8cd932103e6e79625d5f81010b13d1c;
  assign mdsMatrix_41_3 = 255'h4ceb6c296d32909f49626ce1d47e7c4749ac917da89f9570fcc210cd48f9b913;
  assign mdsMatrix_41_4 = 254'h2ca373bdb48253aee65d6cf3167bbb4e69401b30050ace2162b1436c4f1bce24;
  assign mdsMatrix_41_5 = 255'h69b8e20e58d831eaa0c01cc90a049281794320da10f14b0ed68250d9b41b93cd;
  assign mdsMatrix_41_6 = 255'h4f3aa991884f08f08a04ca9f88d8243dc0a04fd6e1afe94780b04356ad6cb7b5;
  assign mdsMatrix_41_7 = 255'h47932258c301bf68831fcc43cc57163b575aff3db144f02aad5d112655471382;
  assign mdsMatrix_41_8 = 254'h34035e2c807c392bf54d603aa4201996df686b0b53e44938ce246b45904c25a4;
  assign mdsMatrix_41_9 = 254'h3127d2106fd860dc5b3f85fbbe8f32926e9509dc614e75f4641a88f5cc88a7e8;
  assign mdsMatrix_41_10 = 254'h2d4b9ebf1e96766f1b919d4f22f4f18c58457de57df091058fbe2010123a350f;
  assign mdsMatrix_41_11 = 254'h2649500e5bd48083bd2e9fae3158d3c9d0c5f70d862e96802e6324c39ce382e6;
  assign mdsMatrix_42_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_42_1 = 253'h1a8baff5dbb13456dbc252d4e5518c1958072609d2948633edfaffc3fecd7d90;
  assign mdsMatrix_42_2 = 254'h25cb8e9a6300f670ecd063ce16b1602d880529ea663e912dce33b7f50212d3da;
  assign mdsMatrix_42_3 = 251'h472b863cb4bb776804fe8b1eb7612a850c6d33eda0ba3c5279fe6cf4ffda4a6;
  assign mdsMatrix_42_4 = 253'h1537a63bb4c7de655013bce70a5400ffb1375014bdfe79ddcaf842a134161306;
  assign mdsMatrix_42_5 = 254'h20e06339136244ff2d99704722a0019ddc00fe04d12eb3e6cc7cf1a1f1a037e6;
  assign mdsMatrix_42_6 = 250'h3f546dc5c7d0ebbe090675f2622513fbeae6c919dd95c295474594e4a0849bc;
  assign mdsMatrix_42_7 = 255'h5f3e518a6e19cda54532b625e43403aeae34c9ef26f7987f39923a84ac2c071a;
  assign mdsMatrix_42_8 = 255'h53f55512feab728ad2cb1dbba78d158feaf9b7b94e3512b3b85ec6d2cc24bd8d;
  assign mdsMatrix_42_9 = 254'h20248b3854c04c6df62dc39500e6c0eeacb9c874afac26c07bd4f1df6fbcf974;
  assign mdsMatrix_42_10 = 253'h1e11ff20c5e78c256e5f35c2bc4455916e9c6a3d31d797e18ef4dcb747ad74fb;
  assign mdsMatrix_42_11 = 255'h731ee02337000c0527225ba0df3648d671e12bb69aba363decd7983d50cb44c8;
  assign mdsMatrix_43_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_43_1 = 253'h12bc354951af77c70eaf1a507868c9d0122797ffa50dbb4135a3c68464c9b979;
  assign mdsMatrix_43_2 = 251'h505d7cf5f3c700b009b92096efe96d88474f2c1018e752b8da793107f9e607d;
  assign mdsMatrix_43_3 = 255'h55c5c57243c224b2b7fe04a06d866b882ee9e91210e7a08fc472eeb13a44408d;
  assign mdsMatrix_43_4 = 255'h55b5a76c9a6279c036c0eb255ac67ef471ad8bca66b5a3e27895b6dd4245ed66;
  assign mdsMatrix_43_5 = 255'h4f3009a64050defcb83cc0cc5109df5c3b3a0922b767b273bd2173147ec00aed;
  assign mdsMatrix_43_6 = 255'h5885965d8fab6a2548c9230ce9766770fb87f1861945b10a924d0740c35475b7;
  assign mdsMatrix_43_7 = 254'h3f9161c38158f00702bca2c4328ba758432f222e114980b13b53367ae58da84c;
  assign mdsMatrix_43_8 = 254'h2646fa73d7b24b95c700a923fecbe6e73e4a651dd9c83eb4f814efae6853cbb9;
  assign mdsMatrix_43_9 = 250'h2c2970094b776854910f703396c62c8b2d9e029c1100a4666e1b29de589bee7;
  assign mdsMatrix_43_10 = 252'hecba50abc6c910c368b5dd3efc2e5075df5a3887d4390407c95595115729581;
  assign mdsMatrix_43_11 = 255'h70843c9b29ab3c80ab270422f3de4a416a4f6fa218a42986a23f93e8859281c7;
  assign mdsMatrix_44_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_44_1 = 255'h51058bc5b5dd259bbd99948277c809b425550f0171dd59ce4e8fcac262e25edf;
  assign mdsMatrix_44_2 = 252'h862d4f06a5805f3317682af39969df9c68d96fd1f0bb9bd633b2a7523f400d1;
  assign mdsMatrix_44_3 = 254'h3f396f261b66eace7fc81087edc967913bac69d3552a2da95365d86b3063515c;
  assign mdsMatrix_44_4 = 254'h3736cfe3d031a1eba4ecbd4e694b6f2102379866d873181252504cd0a95e4c95;
  assign mdsMatrix_44_5 = 253'h1cc6ea7e3e41c7b014148a94ee334aaf7aa65af2ef2f72adc38575610aee0da0;
  assign mdsMatrix_44_6 = 252'hdba801968a54be252f70fe0c9f3649df6d5c6626e34118fd770ff461539fde7;
  assign mdsMatrix_44_7 = 255'h45683db2a4ad0cd63598ca2f9a5bfa5e50701556c864cfce44070f175011365e;
  assign mdsMatrix_44_8 = 254'h24f84477a5a5be1db563f405427fb84699f6a109996c9746294ad2ae8a87fd6e;
  assign mdsMatrix_44_9 = 254'h3622099435b4d99f09e5d0e98877dcea611a9f718fc72cc79e3e241680a0ce9d;
  assign mdsMatrix_44_10 = 255'h52906f9b99251d73f0998e7f58a346890dc5b47e1b27ee4333c15c79e2d7fb02;
  assign mdsMatrix_44_11 = 253'h1141c4c519f83143a2ad47bb07ff16eafa19c8635fe6b70bab4ff0f2b90ceaa6;
  assign mdsMatrix_45_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_45_1 = 255'h5207330378af7d0884eb30da3edd99e2956d5b5fd42214577d919e4a5aa6aadb;
  assign mdsMatrix_45_2 = 255'h6790814fa95bfebe9b1c281166146651a07f97c682dfa115beadbabe7ed729e8;
  assign mdsMatrix_45_3 = 255'h7228f39abd0e7cd670e9cdf51ed4563c62834fafcba8f287c0dce4f59e382fdd;
  assign mdsMatrix_45_4 = 255'h60e94dbb9ee3d6d633321e80fab6f5ef09a227ef52c64940042541cf8df23c6b;
  assign mdsMatrix_45_5 = 254'h3ccd0e88a870900ca48ce21f30b2208a960a17dfd1fdbd8bd92453578d31a4d5;
  assign mdsMatrix_45_6 = 254'h38620584e02567fa7f6271ba39389f57133688399577082d431bc9c5647db3ef;
  assign mdsMatrix_45_7 = 255'h510a094ca7757392addb92bdf9a525975a193ec7e3d0b445e5c0599f4054cba0;
  assign mdsMatrix_45_8 = 253'h139d3abfb2fa8af50805cd042cffd2405cd379db75d313c5b01f7810c49511b3;
  assign mdsMatrix_45_9 = 250'h22ff1dcdfb85ab5560e5205526766b547d31bc3dc40e6994860e07ab511cc76;
  assign mdsMatrix_45_10 = 255'h60c6649176d86c65331ae1380e0ea6d69b5f9f93a89e0a400d48bd936838d452;
  assign mdsMatrix_45_11 = 255'h422be0080d8bc5f063e02e530e8ec025ff981358f26ef1a52926b6da9c97e8a1;
  assign mdsMatrix_46_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_46_1 = 254'h35104dd4683c9da4b8572db9e304394325b7295a3186fd8022207e7306bd7848;
  assign mdsMatrix_46_2 = 253'h1a785a4a959579611ed27d17b3ff5ec62a8c9a5110a9f4a792b67d2d84776580;
  assign mdsMatrix_46_3 = 255'h56745125a0ccf0a806be2375ae07f0083fa43468bcb0f0afacc1289939fa7585;
  assign mdsMatrix_46_4 = 254'h32d1767af64d93f544632964bd1fc368fd651241f1a1775938ad09aaa7362478;
  assign mdsMatrix_46_5 = 255'h4813a7a128a140841216b63238f924ad1c63155efe46511928bb9473c2f7e1b0;
  assign mdsMatrix_46_6 = 255'h4015ade7b07a933a459f700d3287d25d5c1683e0eab6f356362ed38b3063f6c3;
  assign mdsMatrix_46_7 = 255'h69afa60e3c94c934d08f5c39438c9f7bfc1c7bfa01552020ae5e48ac5439bc94;
  assign mdsMatrix_46_8 = 255'h47eca0d0a9a9a404666c93c2a27fb96a73dcc2f64a43befd1d9bf0ea509f5cc8;
  assign mdsMatrix_46_9 = 255'h4eb32afef147f3c1a6ee9d18cd7c16d3a173622607a0a3d674dbe4b76c5d0a6c;
  assign mdsMatrix_46_10 = 253'h1087e38e2848a738a4b2db7e9bf53d1adb19b0c4db6a12dcb0daa1886bab6be0;
  assign mdsMatrix_46_11 = 254'h35f66a96653b73e5ecafdcd414c65dadc2ba87285a332237c2811c809178c118;
  assign mdsMatrix_47_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_47_1 = 252'hd697dccc000a5a96a3d1ada6f2e940199148f107efb770d80b3d25d1599ff77;
  assign mdsMatrix_47_2 = 250'h3dce8da2f81f616deb39ad73efe36f3e4e3836635c2bb8acc1051dcfd48380e;
  assign mdsMatrix_47_3 = 255'h51594257a3cdce7bbdaa362b1afbdff2a78cf11879fb4e5fafde6d81c73e8b2d;
  assign mdsMatrix_47_4 = 252'hf358e63f15702129ed096cb77654473013578fcd1bfddcf8e9e0f23bbe723ef;
  assign mdsMatrix_47_5 = 254'h2e3938aee2b2b375d5d0bf9429489e2d058f1b596c3e401a36093f342ee2e754;
  assign mdsMatrix_47_6 = 255'h5fd3a443602d89c291d0484cd9e05ed7c9ec962cfee029c0de08d086b9f8a28f;
  assign mdsMatrix_47_7 = 255'h65f157b9c895402f5da3f3b52b8f187f2ada31eac1e3a2548aacd09409e1726c;
  assign mdsMatrix_47_8 = 255'h553aa97289b65ca27f30293ca725fb18427113b69a228fc2ad760dfdfac9b659;
  assign mdsMatrix_47_9 = 254'h3d19714265a0b47837920156c16220499fe42b60e3a0028b8cfcd7f967c1132b;
  assign mdsMatrix_47_10 = 255'h63de2442a9b001aca442f5173e7f3e840dd3e0b5c66bd93a1745ffb64e922d1d;
  assign mdsMatrix_47_11 = 255'h72ab9f621b447202c53d5b1128ee53e76da03ebced683a09b5f74f70dd99a58a;
  assign mdsMatrix_48_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_48_1 = 252'hcaec1d4496d6ec4084bcb921343cf4266880d27c73a17e90ac4ad851d0e9024;
  assign mdsMatrix_48_2 = 254'h34c44ca009ffa3843913ee54650d9fd8db1274ffdf9017ec4172f98591bf42a4;
  assign mdsMatrix_48_3 = 255'h472b3d171dc798481820f633bbf949d2de06180417d4844386e6cda5bbed3fc1;
  assign mdsMatrix_48_4 = 254'h36aacb6887db3b9ee0c99b4d9a096f96a9ef3d35bd098fec66d6ae651e2f551e;
  assign mdsMatrix_48_5 = 254'h22d91308111031b76e914a9c32352815700e65326bafd04dc717523c433acefc;
  assign mdsMatrix_48_6 = 255'h5de8ed2ad69749b782972c2d1467ec6e21b5cdb6ec5b8212a9f10c7747a9553f;
  assign mdsMatrix_48_7 = 253'h161f476eee90ce41520bcb80da2200d50553f43ea54e9266e3d6d3cbe4111323;
  assign mdsMatrix_48_8 = 254'h276f86269d259062fa51bae54739408e86f00268298b276307feebf794f9c5f6;
  assign mdsMatrix_48_9 = 254'h2f7af27b015e87639ee0f248a044f683ac5d9cc3f5739306181b5cd1fab37e81;
  assign mdsMatrix_48_10 = 255'h72d993df665d2b5d0f1c186d1156da7d5a494be8af3e95db040bbfdf780f4444;
  assign mdsMatrix_48_11 = 255'h6f9e6bb600cc65992bba0166be23b0a900c773834e2f6b012e18b9e03ee5a2ed;
  assign mdsMatrix_49_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_49_1 = 252'hdfa94d4b9f4156b138d38e34c08f159a1680464d0090a28e7c01a8c268e1e81;
  assign mdsMatrix_49_2 = 255'h44b2deb55408f64b2a336885f4ea04ee621254e8294c2abd337760d1be781701;
  assign mdsMatrix_49_3 = 255'h4c612432d2e684c6b62d3e996ce0279205da26eca770f36d89b5cfd2e7954865;
  assign mdsMatrix_49_4 = 254'h32314750895b8efff12bc528dee5068e7602b333301b5b007e6b2a53c5243ff7;
  assign mdsMatrix_49_5 = 255'h5efc61ea2dc86a54ee5c62cddeecf11c168c260592b58f4e5ad9f611fed22171;
  assign mdsMatrix_49_6 = 253'h11f6b647463593543f99ce3c772fe9cdfcfc76143f3639f034ba9c0f42e84f3e;
  assign mdsMatrix_49_7 = 255'h6421c667c37fd10f182751d25a341d02a8478378e32e3a96d680d2566a4ab104;
  assign mdsMatrix_49_8 = 253'h17c24199dacf47fd751fc024778a1fcfcd21760dcf545a4370668c427921828f;
  assign mdsMatrix_49_9 = 255'h6336ff6e7481cd579a71531d44407ef0fdfcbf5be5118512ef99cdb39c66f642;
  assign mdsMatrix_49_10 = 254'h2c2515841b3af2ba8a0c4a5c4e23b5db67990cf830d5f28b19c790ba97ae40f6;
  assign mdsMatrix_49_11 = 255'h47a15ea3cb7d36ce9a12bccf705defbf47229e720edee6ee728aec3b149eb414;
  assign mdsMatrix_50_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_50_1 = 252'hd2c2b926cf18e52e0ce0f85f63052495c701575d28746a752258e5f90a0a466;
  assign mdsMatrix_50_2 = 255'h411ca94eb7f1336ce8d2322aaca400a19e7c9a68aaca438e18303104e6b5850d;
  assign mdsMatrix_50_3 = 255'h6b25c2fc4068ec9768383c2c6433cb9c09db77450d9b95c5cb766d00bbc2cf56;
  assign mdsMatrix_50_4 = 253'h1942373edb3cab1594347ba87c049f5b63f33c757406c624ac1d95bdbdf9ac4b;
  assign mdsMatrix_50_5 = 254'h23f4f04661a1a48e489a8b0c81a3413b652341ee2ed284747230e945a67b34e7;
  assign mdsMatrix_50_6 = 254'h2fad395bb8540d0fa8f54f1c9234b4baa5fa4e45b5d8931d58005da98826821c;
  assign mdsMatrix_50_7 = 253'h135eba1714c9154258e9655a7a0d560e0073943f4b4715c4e704f88ec20caaf9;
  assign mdsMatrix_50_8 = 255'h6934a94e703a8a0bf9f58d44ff1f7838d80bffb4e5796ae46d043c4af008c6ef;
  assign mdsMatrix_50_9 = 255'h46675d40978cc979dc541ad5c172cd58d72d567a60498e178d6181cca3dbbd01;
  assign mdsMatrix_50_10 = 253'h1d7eaafdcc64996ee3bc1160840efea0ada5909d342b11151d665af8776e6a69;
  assign mdsMatrix_50_11 = 253'h15571811d4c1b1bd96a02caaaa89c49ebd02aba5c04b1b69e60a04c86516c8a7;
  assign mdsMatrix_51_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_51_1 = 255'h52a54019df822918d95159536d6d674ddd1fe3df03464b745d9aab220ba087f5;
  assign mdsMatrix_51_2 = 254'h341c4d9837622e34bc0753e1d96fb6343c5d83cef51039778e201e088aa7a112;
  assign mdsMatrix_51_3 = 255'h66149509b13d680df5ec9871ec7babd0fe411df3d0964612ddce83e9fe1d1e7b;
  assign mdsMatrix_51_4 = 253'h1fdffdd0f855bd02c441b983e36054374e3ca73c1fadcab5026365747910adde;
  assign mdsMatrix_51_5 = 255'h734d4f568af2601d9ea1b0e6471a84f63dd9c48fd3ddea64bad018c07cb56b85;
  assign mdsMatrix_51_6 = 254'h3ce1ed01dd6583122434d7c8d00cc1c82a894617c71aa25c4a847f59e38b73c8;
  assign mdsMatrix_51_7 = 255'h5b71d2a16559ca0827a9694b05aa4bed5da3d7409c26e59842f54e6efe9deb85;
  assign mdsMatrix_51_8 = 253'h1d8dd4935a7bb9a421412f44887cf689b7d9b73aa6e926ed8373ad2257677dd6;
  assign mdsMatrix_51_9 = 254'h2f9fa2e11a72111b4e795980f73e6267f13a14fa42997d6ad4fc73fdef2ccb17;
  assign mdsMatrix_51_10 = 255'h460405af03435caec8f6607895a9647c3a0abbe63b97d659ec935b72178724e0;
  assign mdsMatrix_51_11 = 255'h73d660a1873a2a8da6955cc432471fdb87bb42065dc4ef4beb1f256ad6042667;
  assign mdsMatrix_52_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_52_1 = 255'h5417dfde230d6523b14c5a051a6d0377f2d01a6904ca4781676ade351f7fa665;
  assign mdsMatrix_52_2 = 254'h30eb7de20b951dbac02b56777cdfcde58e421f24f50d2a42c1072883e522ffda;
  assign mdsMatrix_52_3 = 253'h12836f0c09d7ca95339e34164e2ff854b11d8bf3313182aa5baeb85aeeea5d86;
  assign mdsMatrix_52_4 = 254'h3c8d1b41b38e2f4c06a38c6f93cc876901aac63490ce80066b522f8b03ea0e82;
  assign mdsMatrix_52_5 = 254'h3731f088c124267b10ebd8b97e4d201336a78740685e734806b000fcd175718d;
  assign mdsMatrix_52_6 = 254'h291eb5d2a22c696e4e43e626549798ae3548757c3cd6ae78f21fad82ff3b7ff4;
  assign mdsMatrix_52_7 = 254'h284f58e407338b060b8fb7fcdd22afd406788a233c666f67c82edc55ec359ce0;
  assign mdsMatrix_52_8 = 255'h4d14ae81d98e9863238c225087b2501a8819d50d1779f6c41991ca4413ba7930;
  assign mdsMatrix_52_9 = 255'h5b4179657e3f8061b469438ff6dee842fcf1c237a73777737379bb5e1586cf5a;
  assign mdsMatrix_52_10 = 253'h199ebb01ffd2bae9ffc982bcd6b12493dcf05a6c8c005a5be365a3b87f054cb2;
  assign mdsMatrix_52_11 = 255'h552bb44783d6c0962eec52e88eb74d5dea2dd201481da573a2e6f91a8da501fd;
  assign mdsMatrix_53_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_53_1 = 251'h4317f59fe9231a406b3bc83d0be69c62258dc97f1d78dd30c1dbe4c0dae5be0;
  assign mdsMatrix_53_2 = 254'h2f931cd0c56dd755654ee299a1c01956ffe694446a03fc64f3940ecb531b041b;
  assign mdsMatrix_53_3 = 255'h46c916bfc4b8b3cf3ef0bd2d728eea2c18264b25fdcbde725e244e9f8a26aef1;
  assign mdsMatrix_53_4 = 252'hfbfb69cda4e5ebe792e850d27297bdabf001ed24f0e17556abedb279a11a490;
  assign mdsMatrix_53_5 = 255'h5b2fe4b79f97e44f15742ef3f3287533ffd36f0b43621e93a484f33fb1b503a9;
  assign mdsMatrix_53_6 = 254'h260ff72fc1658ad1f7f2d15eca3ad88ba6581e7adb1aefc2b1a8cfced6b3bfdb;
  assign mdsMatrix_53_7 = 255'h59e2ded1f06f61dce4444be315634f65b3fad15cb114349ab0b5b3497ca2d646;
  assign mdsMatrix_53_8 = 255'h5d57d0fbf0c3b8ef76db2bb35c9f493fb25623f649aeb00aac22e1c358719b18;
  assign mdsMatrix_53_9 = 255'h718923fc3ee132fb5fea52feb4290e0e721d67e222691672ceabc383aa018fe5;
  assign mdsMatrix_53_10 = 253'h1cc304a63555e03d85151ec49d65220cce87967e93873ac5538acd062e9bcc94;
  assign mdsMatrix_53_11 = 255'h536748e14c08fb1042074d457c94a032525be9bea9e3cd527dd33e5583706c73;
  assign mdsMatrix_54_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_54_1 = 255'h436c08cf0feba5356afa4aab5302d38fbf4d1fe2169ae4c138cf391f1b55583d;
  assign mdsMatrix_54_2 = 254'h2dbf6e6d0c4b04636c7e660cb3f7c359b0fde1220c3e0d6d4144155362904c5f;
  assign mdsMatrix_54_3 = 255'h46ddafde3208a9cff51ea9751fcb4b6b7f7177214e699b36456673a11787d048;
  assign mdsMatrix_54_4 = 255'h63a9ad375d6ba627f456b47b15b991026d6ad81be48a2d66cac163910cef9027;
  assign mdsMatrix_54_5 = 255'h5f410cb7ea07b5f4d2a48dff74b90b60a9f1cd270e69fd02701ca4e24ec615d2;
  assign mdsMatrix_54_6 = 254'h392453def95a00380dbca6bdf0bfa0cb637d52ba178c468afb588854ba6354d8;
  assign mdsMatrix_54_7 = 254'h3e6556f900cf436cd53ed51bc0778532061f7b652cf3fc4ab9a49e384466a461;
  assign mdsMatrix_54_8 = 253'h18dca3db4c2a346f7621c0270b340b42e44d134f90dd519e5a43112d69b91e94;
  assign mdsMatrix_54_9 = 254'h2ae20616a9981c9f8dd4c5d7289154d7beb3fe11e8f81b41a79fb5100a56f17f;
  assign mdsMatrix_54_10 = 254'h219594e22f14c11ea4d0fb03f6e7f4ad845e0b2b022579061ca5ad4bc55533d3;
  assign mdsMatrix_54_11 = 255'h5a7a8845fb87bcfd91031d0618a489aebe501e6fcc66af764e2411e617733275;
  assign mdsMatrix_55_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_55_1 = 254'h36623261a9ffefce8b055a7550d55b73b9126dc69a54effcb1247db91ef54f9c;
  assign mdsMatrix_55_2 = 255'h4990d842c01dbadb508723adbcca5347d43e891cf177637d7c84d99eaf6c9a8a;
  assign mdsMatrix_55_3 = 255'h64e4ccfe841ca1c735cb300d2b341cd91223eb59d1d4c5397d31f218c7748009;
  assign mdsMatrix_55_4 = 255'h6b389aeb3ad1150e7d47cbe21c8f0eefcada827561d7cbbe16cd032b9e7e85d0;
  assign mdsMatrix_55_5 = 253'h13ad1cc06936aa8398cc74301a956b7954f689e74cad8b6ea6925957387ef8ed;
  assign mdsMatrix_55_6 = 254'h273f33622548fcfb5bf3a2db03a4cb3bd829a5321539a6a7fea65a4210b2ee18;
  assign mdsMatrix_55_7 = 247'h559fa4f1f335846f74a3905f55a80af27c7cf72ac6d4cdea15828c46835188;
  assign mdsMatrix_55_8 = 253'h12d7f1dcda78c6bd345c905e5ea285bcd7f69fa2920157d2be383a6b3b4ccfda;
  assign mdsMatrix_55_9 = 255'h558f3e93ca2b6c1e8c49cecedf197831b23270d63185af35134f88debef8d855;
  assign mdsMatrix_55_10 = 254'h36496379962610698ebce1a63d6181a60eeee0f6ac6b4e21800bb04f87c1688f;
  assign mdsMatrix_55_11 = 252'hde5ae12dd680b5fe058d072062f17d6fce8c64729ff8922e693c5c32286a1bd;
  assign mdsMatrix_56_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_56_1 = 255'h73c1f4fcb7f30104c3c8ffdaa86f27b3f70ed5064f0cdbdd13b13b3f89d89d5e;
  assign mdsMatrix_56_2 = 255'h6d2bf83ec216b78adbb7899ca3a401248948e2ae62b3dfc03de3dcac8ca8cc1e;
  assign mdsMatrix_56_3 = 254'h3a51e31455dc50809e178fc9ade1eef860b8415231e965462492514624924103;
  assign mdsMatrix_56_4 = 254'h3184a52c16a71a87574b65c8699d64850b852010f788cdb124922db124926498;
  assign mdsMatrix_56_5 = 250'h31bf333bfa88fe3caea07f7bede774b13025c000d7d9de200003f4b69692a1e;
  assign mdsMatrix_56_6 = 254'h2e83b4519699fa866c4b532d50c51197a3095f5694edc6f6ffff9a060f0f7509;
  assign mdsMatrix_56_7 = 255'h40570d5616364e81048adc166f1791d5893f15262f9b8f8a1af2f9be6a33dc40;
  assign mdsMatrix_56_8 = 255'h59401e74471fb3190d2698ab7576589a8085e13934b2458d5e507e71a0e49bb6;
  assign mdsMatrix_56_9 = 253'h189769c6567fa7742878efadc204fff5c07786e0b06781e039bebbb56d42bd1a;
  assign mdsMatrix_56_10 = 255'h6c8d0797a943fe3ef3e25ced82a0580866ccfb8c64ac1b6eeead2e155f38c746;
  assign mdsMatrix_56_11 = 248'h888112cc471ab2084f5278e89e6c6cd8ae43865092a629a02d887a77c1bab9;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign tempAddrVec_5 = io_addr_regNext_5;
  assign tempAddrVec_6 = io_addr_regNext_6;
  assign tempAddrVec_7 = io_addr_regNext_7;
  assign tempAddrVec_8 = io_addr_regNext_8;
  assign tempAddrVec_9 = io_addr_regNext_9;
  assign tempAddrVec_10 = io_addr_regNext_10;
  assign tempAddrVec_11 = io_addr_regNext_11;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  assign io_data_5 = _zz_mdsMem_5_port0;
  assign io_data_6 = _zz_mdsMem_6_port0;
  assign io_data_7 = _zz_mdsMem_7_port0;
  assign io_data_8 = _zz_mdsMem_8_port0;
  assign io_data_9 = _zz_mdsMem_9_port0;
  assign io_data_10 = _zz_mdsMem_10_port0;
  assign io_data_11 = _zz_mdsMem_11_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
    io_addr_regNext_5 <= io_addr;
    io_addr_regNext_6 <= io_addr;
    io_addr_regNext_7 <= io_addr;
    io_addr_regNext_8 <= io_addr;
    io_addr_regNext_9 <= io_addr;
    io_addr_regNext_10 <= io_addr;
    io_addr_regNext_11 <= io_addr;
  end


endmodule

module MatrixConstantMem_12 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  input      [5:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  reg        [254:0]  _zz_mdsMem_5_port0;
  reg        [254:0]  _zz_mdsMem_6_port0;
  reg        [254:0]  _zz_mdsMem_7_port0;
  reg        [254:0]  _zz_mdsMem_8_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire                _zz_mdsMem_5_port;
  wire                _zz_io_data_5;
  wire                _zz_mdsMem_6_port;
  wire                _zz_io_data_6;
  wire                _zz_mdsMem_7_port;
  wire                _zz_io_data_7;
  wire                _zz_mdsMem_8_port;
  wire                _zz_io_data_8;
  wire       [254:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [254:0]  mdsMatrix_0_2;
  wire       [254:0]  mdsMatrix_0_3;
  wire       [253:0]  mdsMatrix_0_4;
  wire       [253:0]  mdsMatrix_0_5;
  wire       [253:0]  mdsMatrix_0_6;
  wire       [253:0]  mdsMatrix_0_7;
  wire       [252:0]  mdsMatrix_0_8;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [253:0]  mdsMatrix_1_1;
  wire       [253:0]  mdsMatrix_1_2;
  wire       [252:0]  mdsMatrix_1_3;
  wire       [248:0]  mdsMatrix_1_4;
  wire       [254:0]  mdsMatrix_1_5;
  wire       [254:0]  mdsMatrix_1_6;
  wire       [253:0]  mdsMatrix_1_7;
  wire       [253:0]  mdsMatrix_1_8;
  wire       [254:0]  mdsMatrix_2_0;
  wire       [252:0]  mdsMatrix_2_1;
  wire       [250:0]  mdsMatrix_2_2;
  wire       [254:0]  mdsMatrix_2_3;
  wire       [252:0]  mdsMatrix_2_4;
  wire       [252:0]  mdsMatrix_2_5;
  wire       [254:0]  mdsMatrix_2_6;
  wire       [254:0]  mdsMatrix_2_7;
  wire       [252:0]  mdsMatrix_2_8;
  wire       [254:0]  mdsMatrix_3_0;
  wire       [254:0]  mdsMatrix_3_1;
  wire       [254:0]  mdsMatrix_3_2;
  wire       [254:0]  mdsMatrix_3_3;
  wire       [254:0]  mdsMatrix_3_4;
  wire       [254:0]  mdsMatrix_3_5;
  wire       [253:0]  mdsMatrix_3_6;
  wire       [252:0]  mdsMatrix_3_7;
  wire       [254:0]  mdsMatrix_3_8;
  wire       [254:0]  mdsMatrix_4_0;
  wire       [254:0]  mdsMatrix_4_1;
  wire       [252:0]  mdsMatrix_4_2;
  wire       [253:0]  mdsMatrix_4_3;
  wire       [254:0]  mdsMatrix_4_4;
  wire       [254:0]  mdsMatrix_4_5;
  wire       [254:0]  mdsMatrix_4_6;
  wire       [254:0]  mdsMatrix_4_7;
  wire       [253:0]  mdsMatrix_4_8;
  wire       [254:0]  mdsMatrix_5_0;
  wire       [250:0]  mdsMatrix_5_1;
  wire       [254:0]  mdsMatrix_5_2;
  wire       [249:0]  mdsMatrix_5_3;
  wire       [253:0]  mdsMatrix_5_4;
  wire       [251:0]  mdsMatrix_5_5;
  wire       [250:0]  mdsMatrix_5_6;
  wire       [253:0]  mdsMatrix_5_7;
  wire       [253:0]  mdsMatrix_5_8;
  wire       [254:0]  mdsMatrix_6_0;
  wire       [253:0]  mdsMatrix_6_1;
  wire       [253:0]  mdsMatrix_6_2;
  wire       [251:0]  mdsMatrix_6_3;
  wire       [254:0]  mdsMatrix_6_4;
  wire       [254:0]  mdsMatrix_6_5;
  wire       [254:0]  mdsMatrix_6_6;
  wire       [254:0]  mdsMatrix_6_7;
  wire       [254:0]  mdsMatrix_6_8;
  wire       [254:0]  mdsMatrix_7_0;
  wire       [253:0]  mdsMatrix_7_1;
  wire       [252:0]  mdsMatrix_7_2;
  wire       [254:0]  mdsMatrix_7_3;
  wire       [248:0]  mdsMatrix_7_4;
  wire       [254:0]  mdsMatrix_7_5;
  wire       [254:0]  mdsMatrix_7_6;
  wire       [247:0]  mdsMatrix_7_7;
  wire       [253:0]  mdsMatrix_7_8;
  wire       [254:0]  mdsMatrix_8_0;
  wire       [254:0]  mdsMatrix_8_1;
  wire       [254:0]  mdsMatrix_8_2;
  wire       [254:0]  mdsMatrix_8_3;
  wire       [254:0]  mdsMatrix_8_4;
  wire       [252:0]  mdsMatrix_8_5;
  wire       [250:0]  mdsMatrix_8_6;
  wire       [251:0]  mdsMatrix_8_7;
  wire       [254:0]  mdsMatrix_8_8;
  wire       [254:0]  mdsMatrix_9_0;
  wire       [254:0]  mdsMatrix_9_1;
  wire       [254:0]  mdsMatrix_9_2;
  wire       [254:0]  mdsMatrix_9_3;
  wire       [253:0]  mdsMatrix_9_4;
  wire       [254:0]  mdsMatrix_9_5;
  wire       [251:0]  mdsMatrix_9_6;
  wire       [254:0]  mdsMatrix_9_7;
  wire       [253:0]  mdsMatrix_9_8;
  wire       [254:0]  mdsMatrix_10_0;
  wire       [254:0]  mdsMatrix_10_1;
  wire       [254:0]  mdsMatrix_10_2;
  wire       [252:0]  mdsMatrix_10_3;
  wire       [251:0]  mdsMatrix_10_4;
  wire       [253:0]  mdsMatrix_10_5;
  wire       [251:0]  mdsMatrix_10_6;
  wire       [249:0]  mdsMatrix_10_7;
  wire       [254:0]  mdsMatrix_10_8;
  wire       [254:0]  mdsMatrix_11_0;
  wire       [254:0]  mdsMatrix_11_1;
  wire       [254:0]  mdsMatrix_11_2;
  wire       [253:0]  mdsMatrix_11_3;
  wire       [254:0]  mdsMatrix_11_4;
  wire       [253:0]  mdsMatrix_11_5;
  wire       [254:0]  mdsMatrix_11_6;
  wire       [252:0]  mdsMatrix_11_7;
  wire       [248:0]  mdsMatrix_11_8;
  wire       [254:0]  mdsMatrix_12_0;
  wire       [254:0]  mdsMatrix_12_1;
  wire       [254:0]  mdsMatrix_12_2;
  wire       [253:0]  mdsMatrix_12_3;
  wire       [247:0]  mdsMatrix_12_4;
  wire       [253:0]  mdsMatrix_12_5;
  wire       [253:0]  mdsMatrix_12_6;
  wire       [254:0]  mdsMatrix_12_7;
  wire       [252:0]  mdsMatrix_12_8;
  wire       [254:0]  mdsMatrix_13_0;
  wire       [254:0]  mdsMatrix_13_1;
  wire       [254:0]  mdsMatrix_13_2;
  wire       [252:0]  mdsMatrix_13_3;
  wire       [254:0]  mdsMatrix_13_4;
  wire       [254:0]  mdsMatrix_13_5;
  wire       [254:0]  mdsMatrix_13_6;
  wire       [249:0]  mdsMatrix_13_7;
  wire       [253:0]  mdsMatrix_13_8;
  wire       [254:0]  mdsMatrix_14_0;
  wire       [252:0]  mdsMatrix_14_1;
  wire       [254:0]  mdsMatrix_14_2;
  wire       [254:0]  mdsMatrix_14_3;
  wire       [254:0]  mdsMatrix_14_4;
  wire       [253:0]  mdsMatrix_14_5;
  wire       [254:0]  mdsMatrix_14_6;
  wire       [254:0]  mdsMatrix_14_7;
  wire       [253:0]  mdsMatrix_14_8;
  wire       [254:0]  mdsMatrix_15_0;
  wire       [254:0]  mdsMatrix_15_1;
  wire       [254:0]  mdsMatrix_15_2;
  wire       [252:0]  mdsMatrix_15_3;
  wire       [252:0]  mdsMatrix_15_4;
  wire       [252:0]  mdsMatrix_15_5;
  wire       [254:0]  mdsMatrix_15_6;
  wire       [254:0]  mdsMatrix_15_7;
  wire       [251:0]  mdsMatrix_15_8;
  wire       [254:0]  mdsMatrix_16_0;
  wire       [250:0]  mdsMatrix_16_1;
  wire       [254:0]  mdsMatrix_16_2;
  wire       [250:0]  mdsMatrix_16_3;
  wire       [254:0]  mdsMatrix_16_4;
  wire       [254:0]  mdsMatrix_16_5;
  wire       [250:0]  mdsMatrix_16_6;
  wire       [253:0]  mdsMatrix_16_7;
  wire       [253:0]  mdsMatrix_16_8;
  wire       [254:0]  mdsMatrix_17_0;
  wire       [249:0]  mdsMatrix_17_1;
  wire       [252:0]  mdsMatrix_17_2;
  wire       [254:0]  mdsMatrix_17_3;
  wire       [252:0]  mdsMatrix_17_4;
  wire       [254:0]  mdsMatrix_17_5;
  wire       [251:0]  mdsMatrix_17_6;
  wire       [251:0]  mdsMatrix_17_7;
  wire       [250:0]  mdsMatrix_17_8;
  wire       [254:0]  mdsMatrix_18_0;
  wire       [254:0]  mdsMatrix_18_1;
  wire       [253:0]  mdsMatrix_18_2;
  wire       [254:0]  mdsMatrix_18_3;
  wire       [254:0]  mdsMatrix_18_4;
  wire       [253:0]  mdsMatrix_18_5;
  wire       [252:0]  mdsMatrix_18_6;
  wire       [254:0]  mdsMatrix_18_7;
  wire       [254:0]  mdsMatrix_18_8;
  wire       [254:0]  mdsMatrix_19_0;
  wire       [254:0]  mdsMatrix_19_1;
  wire       [253:0]  mdsMatrix_19_2;
  wire       [253:0]  mdsMatrix_19_3;
  wire       [252:0]  mdsMatrix_19_4;
  wire       [252:0]  mdsMatrix_19_5;
  wire       [254:0]  mdsMatrix_19_6;
  wire       [254:0]  mdsMatrix_19_7;
  wire       [254:0]  mdsMatrix_19_8;
  wire       [254:0]  mdsMatrix_20_0;
  wire       [254:0]  mdsMatrix_20_1;
  wire       [252:0]  mdsMatrix_20_2;
  wire       [252:0]  mdsMatrix_20_3;
  wire       [253:0]  mdsMatrix_20_4;
  wire       [254:0]  mdsMatrix_20_5;
  wire       [252:0]  mdsMatrix_20_6;
  wire       [254:0]  mdsMatrix_20_7;
  wire       [252:0]  mdsMatrix_20_8;
  wire       [254:0]  mdsMatrix_21_0;
  wire       [253:0]  mdsMatrix_21_1;
  wire       [253:0]  mdsMatrix_21_2;
  wire       [253:0]  mdsMatrix_21_3;
  wire       [252:0]  mdsMatrix_21_4;
  wire       [252:0]  mdsMatrix_21_5;
  wire       [253:0]  mdsMatrix_21_6;
  wire       [253:0]  mdsMatrix_21_7;
  wire       [254:0]  mdsMatrix_21_8;
  wire       [254:0]  mdsMatrix_22_0;
  wire       [254:0]  mdsMatrix_22_1;
  wire       [254:0]  mdsMatrix_22_2;
  wire       [253:0]  mdsMatrix_22_3;
  wire       [253:0]  mdsMatrix_22_4;
  wire       [253:0]  mdsMatrix_22_5;
  wire       [254:0]  mdsMatrix_22_6;
  wire       [252:0]  mdsMatrix_22_7;
  wire       [253:0]  mdsMatrix_22_8;
  wire       [254:0]  mdsMatrix_23_0;
  wire       [254:0]  mdsMatrix_23_1;
  wire       [254:0]  mdsMatrix_23_2;
  wire       [254:0]  mdsMatrix_23_3;
  wire       [253:0]  mdsMatrix_23_4;
  wire       [254:0]  mdsMatrix_23_5;
  wire       [253:0]  mdsMatrix_23_6;
  wire       [252:0]  mdsMatrix_23_7;
  wire       [254:0]  mdsMatrix_23_8;
  wire       [254:0]  mdsMatrix_24_0;
  wire       [254:0]  mdsMatrix_24_1;
  wire       [254:0]  mdsMatrix_24_2;
  wire       [253:0]  mdsMatrix_24_3;
  wire       [252:0]  mdsMatrix_24_4;
  wire       [252:0]  mdsMatrix_24_5;
  wire       [253:0]  mdsMatrix_24_6;
  wire       [253:0]  mdsMatrix_24_7;
  wire       [254:0]  mdsMatrix_24_8;
  wire       [254:0]  mdsMatrix_25_0;
  wire       [254:0]  mdsMatrix_25_1;
  wire       [254:0]  mdsMatrix_25_2;
  wire       [253:0]  mdsMatrix_25_3;
  wire       [253:0]  mdsMatrix_25_4;
  wire       [253:0]  mdsMatrix_25_5;
  wire       [253:0]  mdsMatrix_25_6;
  wire       [254:0]  mdsMatrix_25_7;
  wire       [254:0]  mdsMatrix_25_8;
  wire       [254:0]  mdsMatrix_26_0;
  wire       [254:0]  mdsMatrix_26_1;
  wire       [252:0]  mdsMatrix_26_2;
  wire       [250:0]  mdsMatrix_26_3;
  wire       [254:0]  mdsMatrix_26_4;
  wire       [253:0]  mdsMatrix_26_5;
  wire       [253:0]  mdsMatrix_26_6;
  wire       [254:0]  mdsMatrix_26_7;
  wire       [254:0]  mdsMatrix_26_8;
  wire       [254:0]  mdsMatrix_27_0;
  wire       [252:0]  mdsMatrix_27_1;
  wire       [254:0]  mdsMatrix_27_2;
  wire       [254:0]  mdsMatrix_27_3;
  wire       [254:0]  mdsMatrix_27_4;
  wire       [254:0]  mdsMatrix_27_5;
  wire       [253:0]  mdsMatrix_27_6;
  wire       [253:0]  mdsMatrix_27_7;
  wire       [254:0]  mdsMatrix_27_8;
  wire       [254:0]  mdsMatrix_28_0;
  wire       [254:0]  mdsMatrix_28_1;
  wire       [249:0]  mdsMatrix_28_2;
  wire       [254:0]  mdsMatrix_28_3;
  wire       [252:0]  mdsMatrix_28_4;
  wire       [253:0]  mdsMatrix_28_5;
  wire       [254:0]  mdsMatrix_28_6;
  wire       [254:0]  mdsMatrix_28_7;
  wire       [254:0]  mdsMatrix_28_8;
  wire       [254:0]  mdsMatrix_29_0;
  wire       [254:0]  mdsMatrix_29_1;
  wire       [253:0]  mdsMatrix_29_2;
  wire       [254:0]  mdsMatrix_29_3;
  wire       [254:0]  mdsMatrix_29_4;
  wire       [254:0]  mdsMatrix_29_5;
  wire       [254:0]  mdsMatrix_29_6;
  wire       [251:0]  mdsMatrix_29_7;
  wire       [254:0]  mdsMatrix_29_8;
  wire       [254:0]  mdsMatrix_30_0;
  wire       [253:0]  mdsMatrix_30_1;
  wire       [254:0]  mdsMatrix_30_2;
  wire       [254:0]  mdsMatrix_30_3;
  wire       [251:0]  mdsMatrix_30_4;
  wire       [254:0]  mdsMatrix_30_5;
  wire       [254:0]  mdsMatrix_30_6;
  wire       [253:0]  mdsMatrix_30_7;
  wire       [252:0]  mdsMatrix_30_8;
  wire       [254:0]  mdsMatrix_31_0;
  wire       [249:0]  mdsMatrix_31_1;
  wire       [251:0]  mdsMatrix_31_2;
  wire       [253:0]  mdsMatrix_31_3;
  wire       [253:0]  mdsMatrix_31_4;
  wire       [252:0]  mdsMatrix_31_5;
  wire       [254:0]  mdsMatrix_31_6;
  wire       [254:0]  mdsMatrix_31_7;
  wire       [254:0]  mdsMatrix_31_8;
  wire       [254:0]  mdsMatrix_32_0;
  wire       [253:0]  mdsMatrix_32_1;
  wire       [253:0]  mdsMatrix_32_2;
  wire       [253:0]  mdsMatrix_32_3;
  wire       [249:0]  mdsMatrix_32_4;
  wire       [254:0]  mdsMatrix_32_5;
  wire       [253:0]  mdsMatrix_32_6;
  wire       [253:0]  mdsMatrix_32_7;
  wire       [253:0]  mdsMatrix_32_8;
  wire       [254:0]  mdsMatrix_33_0;
  wire       [253:0]  mdsMatrix_33_1;
  wire       [252:0]  mdsMatrix_33_2;
  wire       [253:0]  mdsMatrix_33_3;
  wire       [254:0]  mdsMatrix_33_4;
  wire       [253:0]  mdsMatrix_33_5;
  wire       [250:0]  mdsMatrix_33_6;
  wire       [253:0]  mdsMatrix_33_7;
  wire       [246:0]  mdsMatrix_33_8;
  wire       [254:0]  mdsMatrix_34_0;
  wire       [254:0]  mdsMatrix_34_1;
  wire       [254:0]  mdsMatrix_34_2;
  wire       [253:0]  mdsMatrix_34_3;
  wire       [253:0]  mdsMatrix_34_4;
  wire       [254:0]  mdsMatrix_34_5;
  wire       [249:0]  mdsMatrix_34_6;
  wire       [252:0]  mdsMatrix_34_7;
  wire       [254:0]  mdsMatrix_34_8;
  wire       [254:0]  mdsMatrix_35_0;
  wire       [251:0]  mdsMatrix_35_1;
  wire       [254:0]  mdsMatrix_35_2;
  wire       [251:0]  mdsMatrix_35_3;
  wire       [254:0]  mdsMatrix_35_4;
  wire       [254:0]  mdsMatrix_35_5;
  wire       [254:0]  mdsMatrix_35_6;
  wire       [251:0]  mdsMatrix_35_7;
  wire       [251:0]  mdsMatrix_35_8;
  wire       [254:0]  mdsMatrix_36_0;
  wire       [253:0]  mdsMatrix_36_1;
  wire       [254:0]  mdsMatrix_36_2;
  wire       [253:0]  mdsMatrix_36_3;
  wire       [253:0]  mdsMatrix_36_4;
  wire       [253:0]  mdsMatrix_36_5;
  wire       [250:0]  mdsMatrix_36_6;
  wire       [252:0]  mdsMatrix_36_7;
  wire       [252:0]  mdsMatrix_36_8;
  wire       [254:0]  mdsMatrix_37_0;
  wire       [252:0]  mdsMatrix_37_1;
  wire       [254:0]  mdsMatrix_37_2;
  wire       [253:0]  mdsMatrix_37_3;
  wire       [253:0]  mdsMatrix_37_4;
  wire       [253:0]  mdsMatrix_37_5;
  wire       [254:0]  mdsMatrix_37_6;
  wire       [254:0]  mdsMatrix_37_7;
  wire       [254:0]  mdsMatrix_37_8;
  wire       [254:0]  mdsMatrix_38_0;
  wire       [252:0]  mdsMatrix_38_1;
  wire       [254:0]  mdsMatrix_38_2;
  wire       [254:0]  mdsMatrix_38_3;
  wire       [254:0]  mdsMatrix_38_4;
  wire       [253:0]  mdsMatrix_38_5;
  wire       [252:0]  mdsMatrix_38_6;
  wire       [249:0]  mdsMatrix_38_7;
  wire       [253:0]  mdsMatrix_38_8;
  wire       [254:0]  mdsMatrix_39_0;
  wire       [253:0]  mdsMatrix_39_1;
  wire       [252:0]  mdsMatrix_39_2;
  wire       [254:0]  mdsMatrix_39_3;
  wire       [254:0]  mdsMatrix_39_4;
  wire       [253:0]  mdsMatrix_39_5;
  wire       [251:0]  mdsMatrix_39_6;
  wire       [254:0]  mdsMatrix_39_7;
  wire       [253:0]  mdsMatrix_39_8;
  wire       [254:0]  mdsMatrix_40_0;
  wire       [254:0]  mdsMatrix_40_1;
  wire       [254:0]  mdsMatrix_40_2;
  wire       [252:0]  mdsMatrix_40_3;
  wire       [254:0]  mdsMatrix_40_4;
  wire       [253:0]  mdsMatrix_40_5;
  wire       [254:0]  mdsMatrix_40_6;
  wire       [252:0]  mdsMatrix_40_7;
  wire       [249:0]  mdsMatrix_40_8;
  wire       [254:0]  mdsMatrix_41_0;
  wire       [254:0]  mdsMatrix_41_1;
  wire       [253:0]  mdsMatrix_41_2;
  wire       [254:0]  mdsMatrix_41_3;
  wire       [251:0]  mdsMatrix_41_4;
  wire       [253:0]  mdsMatrix_41_5;
  wire       [254:0]  mdsMatrix_41_6;
  wire       [251:0]  mdsMatrix_41_7;
  wire       [254:0]  mdsMatrix_41_8;
  wire       [254:0]  mdsMatrix_42_0;
  wire       [254:0]  mdsMatrix_42_1;
  wire       [254:0]  mdsMatrix_42_2;
  wire       [253:0]  mdsMatrix_42_3;
  wire       [253:0]  mdsMatrix_42_4;
  wire       [254:0]  mdsMatrix_42_5;
  wire       [253:0]  mdsMatrix_42_6;
  wire       [252:0]  mdsMatrix_42_7;
  wire       [253:0]  mdsMatrix_42_8;
  wire       [254:0]  mdsMatrix_43_0;
  wire       [254:0]  mdsMatrix_43_1;
  wire       [254:0]  mdsMatrix_43_2;
  wire       [254:0]  mdsMatrix_43_3;
  wire       [254:0]  mdsMatrix_43_4;
  wire       [254:0]  mdsMatrix_43_5;
  wire       [251:0]  mdsMatrix_43_6;
  wire       [251:0]  mdsMatrix_43_7;
  wire       [251:0]  mdsMatrix_43_8;
  wire       [254:0]  mdsMatrix_44_0;
  wire       [254:0]  mdsMatrix_44_1;
  wire       [253:0]  mdsMatrix_44_2;
  wire       [254:0]  mdsMatrix_44_3;
  wire       [251:0]  mdsMatrix_44_4;
  wire       [253:0]  mdsMatrix_44_5;
  wire       [253:0]  mdsMatrix_44_6;
  wire       [253:0]  mdsMatrix_44_7;
  wire       [254:0]  mdsMatrix_44_8;
  wire       [254:0]  mdsMatrix_45_0;
  wire       [253:0]  mdsMatrix_45_1;
  wire       [252:0]  mdsMatrix_45_2;
  wire       [253:0]  mdsMatrix_45_3;
  wire       [253:0]  mdsMatrix_45_4;
  wire       [251:0]  mdsMatrix_45_5;
  wire       [253:0]  mdsMatrix_45_6;
  wire       [254:0]  mdsMatrix_45_7;
  wire       [254:0]  mdsMatrix_45_8;
  wire       [254:0]  mdsMatrix_46_0;
  wire       [254:0]  mdsMatrix_46_1;
  wire       [253:0]  mdsMatrix_46_2;
  wire       [254:0]  mdsMatrix_46_3;
  wire       [254:0]  mdsMatrix_46_4;
  wire       [252:0]  mdsMatrix_46_5;
  wire       [253:0]  mdsMatrix_46_6;
  wire       [252:0]  mdsMatrix_46_7;
  wire       [250:0]  mdsMatrix_46_8;
  wire       [254:0]  mdsMatrix_47_0;
  wire       [253:0]  mdsMatrix_47_1;
  wire       [252:0]  mdsMatrix_47_2;
  wire       [254:0]  mdsMatrix_47_3;
  wire       [247:0]  mdsMatrix_47_4;
  wire       [251:0]  mdsMatrix_47_5;
  wire       [254:0]  mdsMatrix_47_6;
  wire       [253:0]  mdsMatrix_47_7;
  wire       [252:0]  mdsMatrix_47_8;
  wire       [254:0]  mdsMatrix_48_0;
  wire       [254:0]  mdsMatrix_48_1;
  wire       [254:0]  mdsMatrix_48_2;
  wire       [253:0]  mdsMatrix_48_3;
  wire       [254:0]  mdsMatrix_48_4;
  wire       [254:0]  mdsMatrix_48_5;
  wire       [253:0]  mdsMatrix_48_6;
  wire       [254:0]  mdsMatrix_48_7;
  wire       [251:0]  mdsMatrix_48_8;
  wire       [254:0]  mdsMatrix_49_0;
  wire       [254:0]  mdsMatrix_49_1;
  wire       [252:0]  mdsMatrix_49_2;
  wire       [253:0]  mdsMatrix_49_3;
  wire       [253:0]  mdsMatrix_49_4;
  wire       [248:0]  mdsMatrix_49_5;
  wire       [251:0]  mdsMatrix_49_6;
  wire       [254:0]  mdsMatrix_49_7;
  wire       [251:0]  mdsMatrix_49_8;
  wire       [254:0]  mdsMatrix_50_0;
  wire       [254:0]  mdsMatrix_50_1;
  wire       [254:0]  mdsMatrix_50_2;
  wire       [250:0]  mdsMatrix_50_3;
  wire       [250:0]  mdsMatrix_50_4;
  wire       [254:0]  mdsMatrix_50_5;
  wire       [254:0]  mdsMatrix_50_6;
  wire       [251:0]  mdsMatrix_50_7;
  wire       [252:0]  mdsMatrix_50_8;
  wire       [254:0]  mdsMatrix_51_0;
  wire       [253:0]  mdsMatrix_51_1;
  wire       [253:0]  mdsMatrix_51_2;
  wire       [254:0]  mdsMatrix_51_3;
  wire       [254:0]  mdsMatrix_51_4;
  wire       [254:0]  mdsMatrix_51_5;
  wire       [253:0]  mdsMatrix_51_6;
  wire       [249:0]  mdsMatrix_51_7;
  wire       [253:0]  mdsMatrix_51_8;
  wire       [254:0]  mdsMatrix_52_0;
  wire       [254:0]  mdsMatrix_52_1;
  wire       [251:0]  mdsMatrix_52_2;
  wire       [252:0]  mdsMatrix_52_3;
  wire       [253:0]  mdsMatrix_52_4;
  wire       [254:0]  mdsMatrix_52_5;
  wire       [253:0]  mdsMatrix_52_6;
  wire       [253:0]  mdsMatrix_52_7;
  wire       [254:0]  mdsMatrix_52_8;
  wire       [254:0]  mdsMatrix_53_0;
  wire       [250:0]  mdsMatrix_53_1;
  wire       [254:0]  mdsMatrix_53_2;
  wire       [254:0]  mdsMatrix_53_3;
  wire       [254:0]  mdsMatrix_53_4;
  wire       [254:0]  mdsMatrix_53_5;
  wire       [254:0]  mdsMatrix_53_6;
  wire       [254:0]  mdsMatrix_53_7;
  wire       [254:0]  mdsMatrix_53_8;
  wire       [254:0]  mdsMatrix_54_0;
  wire       [252:0]  mdsMatrix_54_1;
  wire       [254:0]  mdsMatrix_54_2;
  wire       [251:0]  mdsMatrix_54_3;
  wire       [254:0]  mdsMatrix_54_4;
  wire       [254:0]  mdsMatrix_54_5;
  wire       [254:0]  mdsMatrix_54_6;
  wire       [253:0]  mdsMatrix_54_7;
  wire       [253:0]  mdsMatrix_54_8;
  wire       [254:0]  mdsMatrix_55_0;
  wire       [254:0]  mdsMatrix_55_1;
  wire       [251:0]  mdsMatrix_55_2;
  wire       [252:0]  mdsMatrix_55_3;
  wire       [254:0]  mdsMatrix_55_4;
  wire       [254:0]  mdsMatrix_55_5;
  wire       [254:0]  mdsMatrix_55_6;
  wire       [252:0]  mdsMatrix_55_7;
  wire       [254:0]  mdsMatrix_55_8;
  wire       [254:0]  mdsMatrix_56_0;
  wire       [254:0]  mdsMatrix_56_1;
  wire       [250:0]  mdsMatrix_56_2;
  wire       [252:0]  mdsMatrix_56_3;
  wire       [254:0]  mdsMatrix_56_4;
  wire       [254:0]  mdsMatrix_56_5;
  wire       [253:0]  mdsMatrix_56_6;
  wire       [253:0]  mdsMatrix_56_7;
  wire       [253:0]  mdsMatrix_56_8;
  wire       [5:0]    tempAddrVec_0;
  wire       [5:0]    tempAddrVec_1;
  wire       [5:0]    tempAddrVec_2;
  wire       [5:0]    tempAddrVec_3;
  wire       [5:0]    tempAddrVec_4;
  wire       [5:0]    tempAddrVec_5;
  wire       [5:0]    tempAddrVec_6;
  wire       [5:0]    tempAddrVec_7;
  wire       [5:0]    tempAddrVec_8;
  reg        [5:0]    io_addr_regNext;
  reg        [5:0]    io_addr_regNext_1;
  reg        [5:0]    io_addr_regNext_2;
  reg        [5:0]    io_addr_regNext_3;
  reg        [5:0]    io_addr_regNext_4;
  reg        [5:0]    io_addr_regNext_5;
  reg        [5:0]    io_addr_regNext_6;
  reg        [5:0]    io_addr_regNext_7;
  reg        [5:0]    io_addr_regNext_8;
  reg [254:0] mdsMem_0 [0:56];
  reg [254:0] mdsMem_1 [0:56];
  reg [254:0] mdsMem_2 [0:56];
  reg [254:0] mdsMem_3 [0:56];
  reg [254:0] mdsMem_4 [0:56];
  reg [254:0] mdsMem_5 [0:56];
  reg [254:0] mdsMem_6 [0:56];
  reg [254:0] mdsMem_7 [0:56];
  reg [254:0] mdsMem_8 [0:56];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  assign _zz_io_data_5 = 1'b1;
  assign _zz_io_data_6 = 1'b1;
  assign _zz_io_data_7 = 1'b1;
  assign _zz_io_data_8 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_26_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_26_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_26_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_26_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_26_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_26_mdsMem_5.bin",mdsMem_5);
  end
  always @(posedge clk) begin
    if(_zz_io_data_5) begin
      _zz_mdsMem_5_port0 <= mdsMem_5[tempAddrVec_5];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_26_mdsMem_6.bin",mdsMem_6);
  end
  always @(posedge clk) begin
    if(_zz_io_data_6) begin
      _zz_mdsMem_6_port0 <= mdsMem_6[tempAddrVec_6];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_26_mdsMem_7.bin",mdsMem_7);
  end
  always @(posedge clk) begin
    if(_zz_io_data_7) begin
      _zz_mdsMem_7_port0 <= mdsMem_7[tempAddrVec_7];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_26_mdsMem_8.bin",mdsMem_8);
  end
  always @(posedge clk) begin
    if(_zz_io_data_8) begin
      _zz_mdsMem_8_port0 <= mdsMem_8[tempAddrVec_8];
    end
  end

  assign mdsMatrix_0_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_0_1 = 255'h5903de897b528240d76ed6da10ac7c9f11c7f2705898284780ee4fc16871bebd;
  assign mdsMatrix_0_2 = 255'h635198714306a450cfc8eb9815e3a721f775b5952b232223f0d82966b0d4809a;
  assign mdsMatrix_0_3 = 255'h4d326cfe77392d20a425cea6dda276b78f8fe8ed13ad6aed5151b2c9b1cff31c;
  assign mdsMatrix_0_4 = 254'h341d1346b195b107d0e8e1643db5e9d301511e0365e9d8400103571dcf89f30f;
  assign mdsMatrix_0_5 = 254'h2adf281e9cdf579bdcc2ecf47ffc5947e0cc2ddb3d4648f7080e1ff76d039264;
  assign mdsMatrix_0_6 = 254'h3f9ba93f9112d0adf04613d6ddf4ef276e64627fe2fcc8b974a69b12f14bf5d6;
  assign mdsMatrix_0_7 = 254'h3a56feedceaadefc04e0545a675d9fd5fdcdca99468b0b6d1ff89e13f4439249;
  assign mdsMatrix_0_8 = 253'h1e322952bd57b034bd14fc52bc243684e4698c1fcee6675cbb862911dc913df2;
  assign mdsMatrix_1_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_1_1 = 254'h2d046d99ae08919069dfacfed8d4d756ea4e02e4309c0a34eaeb393ad0ca53e7;
  assign mdsMatrix_1_2 = 254'h2fbc8c14ce0c91d1ec48e4026e34ec7db54de75c08bda96ed7d69c9a0f1ea597;
  assign mdsMatrix_1_3 = 253'h1eaf3f17ebd837f932d47da66c606786b9387f1ee09efdc2cc40e144c8a6d93a;
  assign mdsMatrix_1_4 = 249'h1bb406b1cca87369b0e01136c82f43bbb50eb2426b5aa25358ed8692e625638;
  assign mdsMatrix_1_5 = 255'h41969c6fd623ebeb6d8b9f52967fa0ffdd390c9e24697895908ab68f913b71f8;
  assign mdsMatrix_1_6 = 255'h540ccf5af523caddea704996c6e453167891d23ac871ff9c7f446312fda15097;
  assign mdsMatrix_1_7 = 254'h329584b1c29e31d5a66a9c7eafecf3e460d6e20292d68beabbe36995b3c72edc;
  assign mdsMatrix_1_8 = 254'h353666c2a00f7615111e1efe20f0a0a105f06fa601c59c3cf7f5820c1648ea07;
  assign mdsMatrix_2_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_2_1 = 253'h10db5b64db39b71d6d3ab07616a48af4bf4872dcfa4e2c365beb22d12815875d;
  assign mdsMatrix_2_2 = 251'h6bc4d4ed8cfa94225859d166cd805f67d40f4ee34b2b4ebbb00ac400e5c7379;
  assign mdsMatrix_2_3 = 255'h5be3fc8c1e394698a0d084b00df5f7e38a3bc1d977409b7ee9f235eff4081151;
  assign mdsMatrix_2_4 = 253'h1d749bda31a5aa8f4914dd6652793ca09d32fd2d28e5c5f392ec370eb6b8b97e;
  assign mdsMatrix_2_5 = 253'h1e3c83a86fcf0cd68d6b02db09c3f78da401ff17e6eaca511dc82bb2238f1a7e;
  assign mdsMatrix_2_6 = 255'h6039a5776c4ec52fcd3db6efaed547feccd46962a28d3a409578a9d84b7252d1;
  assign mdsMatrix_2_7 = 255'h48d5ea8ebfc108cea88cacc6ada9cae94147670c9d244d7c93ce65caf2c1a846;
  assign mdsMatrix_2_8 = 253'h169502d77d79521bf65abb2f474cde03ceb3628615614bf902d6bbee5c291db3;
  assign mdsMatrix_3_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_3_1 = 255'h40bc97d4886a5d50551c79a2750c3b30714e30601bfd8b5914c57fa0e03f65a4;
  assign mdsMatrix_3_2 = 255'h67d405857b9ad6b5af87125a1d88ecf020554860df4a87f7712e25ad761a2aa5;
  assign mdsMatrix_3_3 = 255'h6b949fbff1929d6af59f603b840ab48fad5c5105d86135c4f3553551d27d26aa;
  assign mdsMatrix_3_4 = 255'h5fbb4185e67031cbe8aa89e1d9abf4667161ffba883fc2c71c81e52661e1fcc7;
  assign mdsMatrix_3_5 = 255'h6f1ccae7d3513e15cb4ebf12255d0b0317a43bd3886b7c6efdfc9ad5bd85a7e2;
  assign mdsMatrix_3_6 = 254'h38898d282189cb4f84e309b77054cb6124ec32026996898e3d67cdb3853989ed;
  assign mdsMatrix_3_7 = 253'h10ff30ff24f7b525d0e36000756c2d48502c5c9362a8e24c5677bca6603264c1;
  assign mdsMatrix_3_8 = 255'h45d537b3c6b5b23e68a764632ddbfa22dc17e6d70dece753e4746cdf9104c2c5;
  assign mdsMatrix_4_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_4_1 = 255'h6e66ac6db17888cc71115d1407ec75de48c3753ced5f07c4764f7087363a920c;
  assign mdsMatrix_4_2 = 253'h1a8217119c0ba21a6f1edc634d0418bfab5bf3228c3b85e3cc6bd45e2a13f6df;
  assign mdsMatrix_4_3 = 254'h279ef994df8940f7668d3cbbb8f5c49508e21ea3744ba45766ee29c635e069fb;
  assign mdsMatrix_4_4 = 255'h44f0f6830bffed2d42d2f57f701d963674f7d412fd8ce41bc7474a5959fd8a15;
  assign mdsMatrix_4_5 = 255'h6a863955c5636af5d9654ac7127732798e9ba6194ba4b51a6d7da14128e6eef7;
  assign mdsMatrix_4_6 = 255'h4a84344fdf59610c574fc38472dc1f3d1c25c78f0808f98eb641051cfab5ccf5;
  assign mdsMatrix_4_7 = 255'h4c2b28243b35c64e6cbd849b0c2283bc1f1baae5b4b5d4d2e4993335f34ca745;
  assign mdsMatrix_4_8 = 254'h3da0c8c2b59bbc44ff997d84706730350cf1367666fbca2841cea33e03ff3615;
  assign mdsMatrix_5_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_5_1 = 251'h582eefd0d4761f5399f6dfb1018e7338d3dd418276b1fe0236bd49104eb2ab1;
  assign mdsMatrix_5_2 = 255'h71f8fb90f0b91c4c61ff4e217e442fb58ab274627cda765f419ed3db9586af45;
  assign mdsMatrix_5_3 = 250'h32c7f56ad4b73f6517ef3b22dcfafa1837c915c4e88f526a5dd8d87559c507e;
  assign mdsMatrix_5_4 = 254'h3d1691da98244ed018f09e064b951b29bc9bfc79f447d2f81cb3a2f2f2935cd0;
  assign mdsMatrix_5_5 = 252'he8a51d5860eee232eccff3da4c900bf62954f3ee4d76a82e4d3048fe4735139;
  assign mdsMatrix_5_6 = 251'h7de5d39a86deff0767808ff7107d5d6355770877b7d7739092754c837600ac3;
  assign mdsMatrix_5_7 = 254'h2bf50de717e7024842b35cc04ea64622f54b1388e2f67c1fa4612dc2cb49e438;
  assign mdsMatrix_5_8 = 254'h33f51b1afbf182f89a8430b41ca02af8884e39097e5030cb55aaae0ed6de2b47;
  assign mdsMatrix_6_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_6_1 = 254'h25a1c326c17a55c08ec481940e316f5fee035f766f92f7006d80af5a27fae584;
  assign mdsMatrix_6_2 = 254'h22d35a5e070b261c4d94137268f69b6bf9b51202b74435f6b9ade78488d31e90;
  assign mdsMatrix_6_3 = 252'h95fb3bedc09f3aaca4c6feb2736e7813ceda638539fb95fb20b6e9dbabb7673;
  assign mdsMatrix_6_4 = 255'h678c7600f52bb48cbcebddde75edd2949a1bb0276825701430e16fbc88c83938;
  assign mdsMatrix_6_5 = 255'h504d936ab7f0ba0c856a052fbf984f66d9f5db11a1f85d97ddb5af9674928b0e;
  assign mdsMatrix_6_6 = 255'h71bb6f697801bcb9d65e7e6a9d5bd1249d5d48a0088d6af6771827257dfa33f8;
  assign mdsMatrix_6_7 = 255'h53aac0107955449ac949d087a00f9ef316601eae4c3ce5124d37fc00ab3a25ec;
  assign mdsMatrix_6_8 = 255'h649e810f1c3311d8e28c0ed24c9210317f68174dd5471455d4b976d085da3a97;
  assign mdsMatrix_7_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_7_1 = 254'h291e973dd6aa457eaf1ab8fda9c2ca1f902baca3610da95ea2eeb45a393b5d61;
  assign mdsMatrix_7_2 = 253'h19f8db696f217293d3602c1bd341acaa71718572953a4f31534144b3127ecf50;
  assign mdsMatrix_7_3 = 255'h5ae0fb3df61c0403585f8808b5f370fd38a91b0bb4e04e0d8b489166a9f7fda7;
  assign mdsMatrix_7_4 = 249'h16de3ca6fe0fedde3ed1a2e372435be5bcc597f086c3fe095fa129b41c08583;
  assign mdsMatrix_7_5 = 255'h57397ddfad5fcc05f42214004eab3e961f39f95be97904665644b8a20e40a015;
  assign mdsMatrix_7_6 = 255'h70072fcb20784dccc318b93cd7c6a5ac4f208e94146b27140bb3188780978da1;
  assign mdsMatrix_7_7 = 248'hae2e451071caf6da89f20f1f13770fd1652ff49704e9dd58a18a0d30b87add;
  assign mdsMatrix_7_8 = 254'h3db23e80660e70965ba3251292c5d0465fb4c0c8a074fa4fc5fa146015602b37;
  assign mdsMatrix_8_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_8_1 = 255'h48beaaa5e89e3954fc404ad809a60dd5a31667486d86b2d2544cb86ca72f8008;
  assign mdsMatrix_8_2 = 255'h547d286ca911913daa90421ac2502a39a372cb9f660c86960c64c8e909b8b0df;
  assign mdsMatrix_8_3 = 255'h6a0f6499f1ec2bf5b871f693469ee3cbba69e0611ea368c1fd66bc07ed510cfa;
  assign mdsMatrix_8_4 = 255'h44666c0b0b8934fbfbe676b470e13fb8edb5bbb53c5cef7e5abec89e40965878;
  assign mdsMatrix_8_5 = 253'h1b3a81625455c49ad5fc858f868330556bdb6d57293d4803e5fd0d15b86f27ba;
  assign mdsMatrix_8_6 = 251'h53b0a68a79ee10131be74877f78414513199e66b4debd35cf5e488d3607f523;
  assign mdsMatrix_8_7 = 252'hdede8a1ac2fa9293a67d42b749bd7da701d697d354d3897163f728d48df85bc;
  assign mdsMatrix_8_8 = 255'h6f8e98ce827eaa57a9aecd78b667b38c168d9ae51ecd7e9bf919e4836eaef484;
  assign mdsMatrix_9_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_9_1 = 255'h6da8b4065138e7192679f939a9f1e32a250b08294f1cc08c21e82f1453420859;
  assign mdsMatrix_9_2 = 255'h5c2eaeb071fd1ab18bffba9f05e1c2576a1644b8abe9db6477b0045cb8b491cb;
  assign mdsMatrix_9_3 = 255'h4c46b27ff0da12934dc5414531cb56dc1966062179bf9f68468b5b7bd227784a;
  assign mdsMatrix_9_4 = 254'h25d2d5baefe640820acfbc6570340502ae75e87ae6c6f64201ec12860fd94a74;
  assign mdsMatrix_9_5 = 255'h63940a6494a785168e4957a86a0c80dc0becf343a26c381fee2b8cd9f5095138;
  assign mdsMatrix_9_6 = 252'h85b88413cfeddcc34c727d697b4546f5351c4b02effd1af894f17d9bd46c2ad;
  assign mdsMatrix_9_7 = 255'h44d953a272039d7fe57af646f2ef125dae5afb1a9d1fafe098ee58adefadb056;
  assign mdsMatrix_9_8 = 254'h3eb37ceb1e53e7e208b25bc03ac70e460c74b56c8ef8ed6ab670052d7633352e;
  assign mdsMatrix_10_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_10_1 = 255'h4551420a7bbfb7808282a907b23059d19e806bb73a6fac989526c1b8b1c58c1f;
  assign mdsMatrix_10_2 = 255'h6e4c8eff2dde690557dca18aa8cce810e300cd524ce4129b78fef45995d37d0b;
  assign mdsMatrix_10_3 = 253'h1aaff22170ff74267668cf831a010898e6faffd0d9a33a0279f8db0c354b5a18;
  assign mdsMatrix_10_4 = 252'hb0b667f84eb4bddc853cc7cd7b02c799e1dd4a7865ecffd1e7f1d2e5a4ae951;
  assign mdsMatrix_10_5 = 254'h2d141e1fe923fdafc586d9e4fddf00e53a1b3541c998e5ba64baa37b894e7392;
  assign mdsMatrix_10_6 = 252'hcffec28f5e221e815ab8b6c7cd0c56a66c4f43f8864ce2f2e652dd038f718a8;
  assign mdsMatrix_10_7 = 250'h216cf757f4b94f5e46bd7bc9be628522f7ed7b07bcbc92dc82201ebd261399a;
  assign mdsMatrix_10_8 = 255'h620b1d3c48c36f0df34d667b0b72ea91a9ca78c713c42f774f8f95ef249a6666;
  assign mdsMatrix_11_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_11_1 = 255'h6594fd15ff2b1a1e92c5d3188735424b714e646a079cc44f441b8b4b547546b1;
  assign mdsMatrix_11_2 = 255'h4c8d4399560c1e73bef09fb16d78803f03397cb852da11d6037cc83f04f5acd2;
  assign mdsMatrix_11_3 = 254'h3ebb585b4203e35bce7de42e268f585dd1c683e0b9c11239174dc9e0cd5a449b;
  assign mdsMatrix_11_4 = 255'h71f4d8fbf7d9ce82cfff055b72d61b3e19ccfd278fcab736a37f0aba67015731;
  assign mdsMatrix_11_5 = 254'h2647f7f0e47f6f0fa00bd1c4a3196fb3100d6863468fc5ca8df3d14a03261fc5;
  assign mdsMatrix_11_6 = 255'h6f012b71ea9f15203db73168e95f026226d771bec90e3e8b4c955574852f937b;
  assign mdsMatrix_11_7 = 253'h11bde248b75b5e3afe82b9eb5b96abdd896cc2f96a21ec8a4ac1f3f641c4e188;
  assign mdsMatrix_11_8 = 249'h1903bb4dbab74d3d382412fb5316e71483a1b10235460637d04e731a85f146d;
  assign mdsMatrix_12_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_12_1 = 255'h7108dcdbf70710fa8fb338d2e5b5631f26ff652c62440a457cb8fec168c91ff6;
  assign mdsMatrix_12_2 = 255'h6e9fe2d4c11f23c1c31a8d61b0a6f10cfa34d5559099f10e49ec494090f343c2;
  assign mdsMatrix_12_3 = 254'h2c3b4ee7c7d23158a00040cece9e79ffaf4e1a4e236ffefdb7ed75762e958069;
  assign mdsMatrix_12_4 = 248'hc566527d4113ffd55a415febba92baae0d6bc3224ab139bf0f7989c6517d9f;
  assign mdsMatrix_12_5 = 254'h3dc3d2318330ec1403c85de6349f8bdc9a9363d9daf420f3d423f87f61f6f7d6;
  assign mdsMatrix_12_6 = 254'h348d4c505e82177ca1d1cc001a881b5ece76f5e5ce2c45cde699d3bd41a64dd7;
  assign mdsMatrix_12_7 = 255'h4bbd2a709c57149ea88acbcad9cb6929f5586f15aed76f3fc8934e9b891f8247;
  assign mdsMatrix_12_8 = 253'h14cfcbf06ece9cb0b852c58753374aaae83aa4dbc5f7178c95ffdc1f61122406;
  assign mdsMatrix_13_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_13_1 = 255'h53f460377eee398ceeffbdf8913610a2a2d8bdf45d96c28045ed22e26313569b;
  assign mdsMatrix_13_2 = 255'h717a123b2f3652d24f5390f5b058b7787a340ae227584e22b64e56e3f9ac8f2c;
  assign mdsMatrix_13_3 = 253'h1925583d3aa55af369d9923327ffca04cd99e138463f2988cd372e9b4a757af6;
  assign mdsMatrix_13_4 = 255'h725755cf65b20b1f5a8f8500efdce262ee1bffbf902ebf84f7aadeb14f5074ff;
  assign mdsMatrix_13_5 = 255'h45f0196161f5cb16609cee58a7c1564ce0af3403c40cef7f75e3483f758429e2;
  assign mdsMatrix_13_6 = 255'h50a786296c33a3d82b51fb59516781937f37bc40a3b6f1fa8609a987bdfd0662;
  assign mdsMatrix_13_7 = 250'h218bb54576393573dcfafb33d1673f8c94d3b1072d376a0aeeb3025ff00ecea;
  assign mdsMatrix_13_8 = 254'h3be2538f94b3a18703182ec587bb150a7b60f75a654909593d8b8de1e38e9b0e;
  assign mdsMatrix_14_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_14_1 = 253'h13174fabcf54231268b458eea8d03d63b8b8e4a255308981baab93768db4401b;
  assign mdsMatrix_14_2 = 255'h446251b75f7cf8b7633794fca16f176e4a254aeca1847fc950e3e8b7605c6024;
  assign mdsMatrix_14_3 = 255'h6de125c60596e620a28c84eecdb9a74fddb47821be6141ec7f00b2cfcf225915;
  assign mdsMatrix_14_4 = 255'h52f69a8c5d67ff5df093d109db731ee70416c85c21181f7da7a7ca54092010aa;
  assign mdsMatrix_14_5 = 254'h2e05e7b3188f95eb7722d03f3205b641216c793cc1d7fd7a0f2e72c139a0418f;
  assign mdsMatrix_14_6 = 255'h6ba49194797db52d62c0a56e686e4341a21d3966a3e3e1c1fb8c654bc4499b60;
  assign mdsMatrix_14_7 = 255'h736933a7ca0fff4cc0412e2ec35b7d4149a0ad7df7a11026c35610f0a7ba7fad;
  assign mdsMatrix_14_8 = 254'h27b8992db5a48b4715d7dfeb489ed9b367a5c4043a26654ea6a3a98d5cdf722a;
  assign mdsMatrix_15_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_15_1 = 255'h5802a391ac1262861f22d5b4305ca61bf39182fe6becc1352862918246052f2c;
  assign mdsMatrix_15_2 = 255'h5e660ad0c6afe3cb798c4773037acce4ee5355c767b4249c9f839db985e9f084;
  assign mdsMatrix_15_3 = 253'h1fcecb086b5a022aaa1b55014e2331f503e63fea388a2775e73c02be23a09d90;
  assign mdsMatrix_15_4 = 253'h1ad72d2cf2009a59af514e8315c4b82b37f209b786c5d9277e34564c6b004908;
  assign mdsMatrix_15_5 = 253'h1d6ce64319d05a6753143de2e8c98527aae3d08ae9736661d4d44a30a54deea8;
  assign mdsMatrix_15_6 = 255'h455ad7b42f4406107eb1c0a63ad56e5973cdbb4a237f3c513d38a06ed9eeadad;
  assign mdsMatrix_15_7 = 255'h70216cef87b0328d3f70d4f984ea9610eeb3322b208b572c1d66a404edcc6adc;
  assign mdsMatrix_15_8 = 252'h82cfdee3e2a71cc8f07bda119e7c41de9c28b34aa3358ee4750fe7352a710a9;
  assign mdsMatrix_16_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_16_1 = 251'h729e491e4970589de51c7dba33cb7481923c595e33731eeaab68c43d2997498;
  assign mdsMatrix_16_2 = 255'h6c6223def3cb13a0e9b644e76cebac5c1c1b6a28fcdfe70d35ce0864af3d1862;
  assign mdsMatrix_16_3 = 251'h7173e3a97206681df8d827d4885888de29ea75f41aa84fb39812fb0067a7137;
  assign mdsMatrix_16_4 = 255'h5932e83fe09729a5ac9ba64b0a444352ac51a2d0d2590aac4dc6208bc8a0c1c0;
  assign mdsMatrix_16_5 = 255'h49cf9968f73791fc7d686e76ab75f661da68791883603655030d66128ebd5368;
  assign mdsMatrix_16_6 = 251'h6c92d778523d7ba97b30836ef6d7acfba598963d036eb64b44bf9757a0f22ed;
  assign mdsMatrix_16_7 = 254'h3529ea8e60780fd2e9c088d205075fe64e60623e50fec058586e9fcc5e1d8823;
  assign mdsMatrix_16_8 = 254'h39ee14d5403dbbbacee1033ba037258c50f9606cc9758df787db93b4144fb62a;
  assign mdsMatrix_17_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_17_1 = 250'h3c433330469ebd8194e56a7a7d9b4c95cebc81415ce7ae1c39096eec31e6c4b;
  assign mdsMatrix_17_2 = 253'h1134d998e7e84bb2a8d65bbbe7101e2b0295f289236cfee4aa5403df32cf6d18;
  assign mdsMatrix_17_3 = 255'h4484f625a450d3ef59f4f415972540fc5418264a02f3d4a0539edca318543a28;
  assign mdsMatrix_17_4 = 253'h15d7e14d1b6c457dc4917fcab89ef6a244c79f6be7aa47d63f348ad470da5e11;
  assign mdsMatrix_17_5 = 255'h6d4ae3db01ae57412ca3d05b396383f70aa0dc2359a4b13328f8e459d74a96ed;
  assign mdsMatrix_17_6 = 252'hb2a9e006ca1eae4dce2dbf14aa672c56d29d6ebe1a77028811cf46f0afa1b24;
  assign mdsMatrix_17_7 = 252'hbebb1e1bdc2eb121551d50fe99867d28de245d3f304a0eedf4af1ec44eafc60;
  assign mdsMatrix_17_8 = 251'h745ce27b7cd49a589d94c89041cc187f8a94e96cd7210a9b5062b45a577d394;
  assign mdsMatrix_18_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_18_1 = 255'h5bfdd066d41ffa32f264eebefb6cd4c1fe98f347182ebf5613984baec066fcb8;
  assign mdsMatrix_18_2 = 254'h253992fe728ce4e987009b0487a436436e5c7b91d302352eceb060e583ef4f8e;
  assign mdsMatrix_18_3 = 255'h5b404017068fe3f8a1c464109606599f91553639ce1ef0f710da863e45951845;
  assign mdsMatrix_18_4 = 255'h6f9006e477f387303bbaa26a645d54c6328d28819c5183d8457159a1b09aa2c5;
  assign mdsMatrix_18_5 = 254'h333097f70a44738d5d8f872b610cfbb4599225d4935c7f574b5a044b98307845;
  assign mdsMatrix_18_6 = 253'h154193ad6649ce1377fffbc7aef9abd830f9847ff4a6159060a855c9498b1947;
  assign mdsMatrix_18_7 = 255'h438ed1ee3e9c0974032b056353b07b6efa66f36fad9774f23b3adab133937858;
  assign mdsMatrix_18_8 = 255'h4536fee7f6be42664f671bf48f0a0fb902d5827371e30f3ae4034e4a0756ca75;
  assign mdsMatrix_19_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_19_1 = 255'h53d31871f941a70a6f6b4e80e93ef2160a2f7c47259fb643827f8afdb1f548db;
  assign mdsMatrix_19_2 = 254'h209aaab4636cda28bf74444fa5d94c71454b101a362049c30b71c5ba5c14b246;
  assign mdsMatrix_19_3 = 254'h3d1bfd7e0d7def0398f2239f0947d00a157edcf417c6e64e87551a55edf860b4;
  assign mdsMatrix_19_4 = 253'h1499c8ad19f02b07543a10040b9db2458b1f39a41376e7239006cae73ba43e68;
  assign mdsMatrix_19_5 = 253'h17da918b381c252efcc6bc1a4a1f28a3f8cd1a13d90170ab40a61b6fc042abbe;
  assign mdsMatrix_19_6 = 255'h5b79087d4850d71d02823e1236a5d10b8bb67dc07e90cb16de27f0b294842886;
  assign mdsMatrix_19_7 = 255'h6b185803867e116ea33d4e9ca0273b5e8a638acc3b8128a40f5ee618d69fa8eb;
  assign mdsMatrix_19_8 = 255'h5eb03931c76b405e972b5b23ce3518a0e470bd03561278e3fd3d6a5591751828;
  assign mdsMatrix_20_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_20_1 = 255'h70fb3f1e74ec97d278767f72a54d7f7bec9e88fc075dcc775e4fc4a2399926de;
  assign mdsMatrix_20_2 = 253'h1048eb0ff0ceafab229dd18020314f231035d8cd0146239ceeba9a29cc4aac6d;
  assign mdsMatrix_20_3 = 253'h14225b34bc852c147138c8bd01525f66e4d9dc9172fe680994f8375cf62453df;
  assign mdsMatrix_20_4 = 254'h2ce478e57211d8216b154282705e8b9e0b646b4d0a180eeb0ed790b2f52af609;
  assign mdsMatrix_20_5 = 255'h474d8f38894f21fa168323d5b5d6f19c59f5cee438f1567d5ae9bb02d5669896;
  assign mdsMatrix_20_6 = 253'h10502b3c97a0ff7cb80541863025de4ba5356f920305ba639d70a91296a25061;
  assign mdsMatrix_20_7 = 255'h5beaeae3bf71a7eaec2f0cae18d420e8fd27b2dc804c1487da39fe5023b8198d;
  assign mdsMatrix_20_8 = 253'h16ba28fba8046811ae5ac8e72b440cb922757924240a9bd0ff71ffd51a100bca;
  assign mdsMatrix_21_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_21_1 = 254'h2f13e16e93824c3937c5c82e3b44047b8d77e498d7847e0965ada90d546eb468;
  assign mdsMatrix_21_2 = 254'h3fbc2035575203ed23310092ac78fd9874561935a66f253496409d26985016ff;
  assign mdsMatrix_21_3 = 254'h3724e7f345a7a2a38cca26e89c8fe3a908f0a77683078c3c21913598a7b620dc;
  assign mdsMatrix_21_4 = 253'h1f20e79f377d1fea86caf84564ddd129e16c7897e8f5accb213dc7e6c3b584bb;
  assign mdsMatrix_21_5 = 253'h1f5e502e47c87fb0ea7e8eb8c9cc404cb24b42b299a75084f207ad63b352330e;
  assign mdsMatrix_21_6 = 254'h3065a19ef5cd37c00ac27f8698aa5160d00edc9fdd35a516e96d0695f2d26363;
  assign mdsMatrix_21_7 = 254'h271274ef65972da4b7af13eca79b7ed5039693a0afe39e34e2ee0816f933d545;
  assign mdsMatrix_21_8 = 255'h402bcea8a4ffe961e4f527be070a8700af31b4c2c73edf1c11122c98d7d2b3a9;
  assign mdsMatrix_22_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_22_1 = 255'h67d6fb4c34a3c4dd342295d2ec64729d76499d1d4d359a369f8f4a63f0ead220;
  assign mdsMatrix_22_2 = 255'h64a7fd10285d477a041d70fabf9180cfbbcfb310a783c3b7c2f4de4c859c7a3a;
  assign mdsMatrix_22_3 = 254'h23c7410e23b75543e4301ada27cc3f45a6e363617aea156df56e3cfaccdf594f;
  assign mdsMatrix_22_4 = 254'h396978323f2ea7849d1c27892ca2de8c6d47a519669d1bf5d0042efa56986d0d;
  assign mdsMatrix_22_5 = 254'h3b791a044e4652053a45392b50fb2ea670f8a4cca6933e04225b6033f03c8483;
  assign mdsMatrix_22_6 = 255'h7039581f5209af41ef569b991a5e358ed704d66d1d3365fefa7a50fd017228de;
  assign mdsMatrix_22_7 = 253'h1ed0e13ab872789c585040725a4df4547e58312e802bd7b990910f5397a5cb8d;
  assign mdsMatrix_22_8 = 254'h3e13ac7e05adc1ae00ff6f796d810f6920f6015f1d65b4cf56ba91bb04d35fcb;
  assign mdsMatrix_23_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_23_1 = 255'h4f59578f940154c10b2a7508ecd4fb7979b8786bf59d4a01df01a2a5274d0725;
  assign mdsMatrix_23_2 = 255'h5e0e2dbb43667db9be569e3eac3e35b99bf09a4819b2c53518ea7ec315d1d79a;
  assign mdsMatrix_23_3 = 255'h536ce77acf6dda3a310ef8aabedcf16432deb58cd7d942da5c9abc77e6aa11c5;
  assign mdsMatrix_23_4 = 254'h3b3c02f28f6e79c451a187e628d6c36c8a5e9070cb52d482fc1c3d5dd87e7735;
  assign mdsMatrix_23_5 = 255'h642b01172dcbe45b400de5c2a153185a12892104cb3274b22f87a95e005fc331;
  assign mdsMatrix_23_6 = 254'h2e6015f148784ecceb1674aabe06b5d9e0dd0d0276c490eec8b6e9d6a26d8c05;
  assign mdsMatrix_23_7 = 253'h102669d4a1a08e0ea4cbf891dbf5c488f4eaee8c8bac5aca29dbf74d94be0305;
  assign mdsMatrix_23_8 = 255'h6ff516c93ac4fd2e20d6a01d60c3740b0c0c123f9a44c585158a84bc5a52f637;
  assign mdsMatrix_24_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_24_1 = 255'h538a089b30064f61e277afa77f04273a52e8edd30a7c0a879748c33ccc5b7249;
  assign mdsMatrix_24_2 = 255'h4870af813f24b3c8d2987e519e9ad62f01addddfa4dcf1e444a248399ea20711;
  assign mdsMatrix_24_3 = 254'h3315267e1415930fd1a581e79d95d948a894ddfe7ced0bf038ac80f03865afea;
  assign mdsMatrix_24_4 = 253'h190b0bf48b85e061ea59f3781a09733265dfd007469dba5807d724aedb14c1d4;
  assign mdsMatrix_24_5 = 253'h16c38935a542c9dbae0543d20ede5a545f8511321de430634eb53e25f831092e;
  assign mdsMatrix_24_6 = 254'h3c6895762dbfa5ed53ddeb5e788aabbfd2f994ede84187c0eab559d6318cf543;
  assign mdsMatrix_24_7 = 254'h3afef7c4279ec9433f346e5c565ed75da6d3e548d074e617c087407e58f96d2b;
  assign mdsMatrix_24_8 = 255'h4105ba46416568d865c1b21efc897d1276a655cbcca8f37c747bcee6503529a2;
  assign mdsMatrix_25_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_25_1 = 255'h6ab5102bee7e8c1fd8f29420d005b500fdaf27e3b7e468e1cd5a8432025e1bf6;
  assign mdsMatrix_25_2 = 255'h614a2f98e04e1d1483978ce8b1501936d49d6e22f426fb3f5408dd848ad30f90;
  assign mdsMatrix_25_3 = 254'h3bedbd669d9c0de5cb901988375348084a76107940822d1260b2f5dcf26a7897;
  assign mdsMatrix_25_4 = 254'h3a2c733385e3330286f1c85a9bf4769175a02c0aa793c914a923ac0b0568d008;
  assign mdsMatrix_25_5 = 254'h33171c56f4fdccb75b8d3fa03fbe14b3ac32ed424069f22c7191037de2dcb94f;
  assign mdsMatrix_25_6 = 254'h253b993a3983c9a1a0a588a1ac1771f4da994941527536503a2bdc29351514d1;
  assign mdsMatrix_25_7 = 255'h48dbbfbd9184df28d20d0726e452b1e739d401400bca995000672dd84ca68fa0;
  assign mdsMatrix_25_8 = 255'h5132edf61108340624fea82ccd9d813b9eeba3497de005c681597b7d6c974a5b;
  assign mdsMatrix_26_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_26_1 = 255'h673b35557053cb4c9b12d31e95ad55668b60e6e648e2a64f1ca5a4a13e16f86e;
  assign mdsMatrix_26_2 = 253'h1a979ed2aa3ab68c953d07bb82d0ea6df707852288501ad43761f72954a79cd6;
  assign mdsMatrix_26_3 = 251'h7601d0b2c0061047c6ad63a2d691569109616265fe016885f81af472cb54f44;
  assign mdsMatrix_26_4 = 255'h4bec09ec76d421eba53539b556f13ca16125f1fb045eac36bfc16d7e3478ed0c;
  assign mdsMatrix_26_5 = 254'h262895efa8214a2ddae45906147a7ff2fc001870c3187f17ee4f518b59adb0bf;
  assign mdsMatrix_26_6 = 254'h3532841c0cb28cc2a06c420f55f703513e6ce39f52bb1acfbae1e18bd80b5f73;
  assign mdsMatrix_26_7 = 255'h4a52b675bda4e0e0c025d5dbaa61dcc1b2263899ced7c31d7db4c960467efd52;
  assign mdsMatrix_26_8 = 255'h54fbd039c37d5991f1c468c93b39a80e35980e4789180b6f7eb3dcaff299df3a;
  assign mdsMatrix_27_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_27_1 = 253'h1df327c1b5b7ae333724f3f9010d80b274ad4dd6db0d5bc377e962a9923fbe97;
  assign mdsMatrix_27_2 = 255'h54178e493ccac4d6e5e75b1154b671e6698e2692fb30b3a0f563e4f8e13bba44;
  assign mdsMatrix_27_3 = 255'h6fcffcc02a10ce8fb3ef47b43d180c37f91ddf97ef0b0c3d9657bf6d064576c0;
  assign mdsMatrix_27_4 = 255'h492954e815ff3cfd4299b9f6418183f164cf44e287de51b152cc2ed410f96bf0;
  assign mdsMatrix_27_5 = 255'h4566ebc22b24491d59f9b5a393e23745074dbc7dbef1323210faff9450d76f49;
  assign mdsMatrix_27_6 = 254'h3cec81e23ba89725dfee926015e9ac0fd48399855c590b879af01ccbb219a8fa;
  assign mdsMatrix_27_7 = 254'h3dfc7e1cce63b3db741d069b0ab3783bbc63a69c71623599934dfd0ce0ebb26a;
  assign mdsMatrix_27_8 = 255'h587a3d67116f13efe786e2bfd5cd9a32c21c3550d63243cb0a4a241bc7568e05;
  assign mdsMatrix_28_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_28_1 = 255'h6bdc170632586211dd440c3568bca65828591a2e02464d601854edc6b6ef7d5c;
  assign mdsMatrix_28_2 = 250'h2cde2f349c9a3dee569bf7ff9ca652dc01cada820b7fec4b56efb824d562485;
  assign mdsMatrix_28_3 = 255'h508fb93494fdb29f043da38fba427d4610264f9f00d47458bb410424bbeef003;
  assign mdsMatrix_28_4 = 253'h13e1d80335d7a54963900fc460395574df830e01cba8fb81a9f7bf34525231ee;
  assign mdsMatrix_28_5 = 254'h206c6e7f739fdcb5d63f61256fb820a0ecb83230bbff440f44d784a70ebdf659;
  assign mdsMatrix_28_6 = 255'h5fc14b842e7b40bbef7033bd433972544a752fdce97d6bf65cc160cc02f769d4;
  assign mdsMatrix_28_7 = 255'h4c7924f2e6426a3d73536a6e2cdad6cec05f215cdffb238e837c39891f26267b;
  assign mdsMatrix_28_8 = 255'h5a75b1a52617c509f5a43ba408a8290eb984336a82167ed8d69c9ba56eced9a4;
  assign mdsMatrix_29_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_29_1 = 255'h46014a6f9de92a1add7f0781dd24d267aeb7cb229c6c0c641f6047e025c02b54;
  assign mdsMatrix_29_2 = 254'h2cdc2d174ad36971f2478347a696c389fa6b07fdcb4ce121f1e893907e702072;
  assign mdsMatrix_29_3 = 255'h539b129a641a4ffcdd69e0c76ab4b6bef2c72cc4d05d17dd4d79da55417d710d;
  assign mdsMatrix_29_4 = 255'h53ee52dd3d57d260e2d281b902527c19b79a93e5e084c2453684ba39344a5a8b;
  assign mdsMatrix_29_5 = 255'h415b25e34a8773a383c6d68bc978749dc8828ffc1fb61a17375718935cb79dba;
  assign mdsMatrix_29_6 = 255'h422a19718833ce216357df947688cc5bcb2d7b3edb67e4434b9f8f04a4995d55;
  assign mdsMatrix_29_7 = 252'hc41adcf6ced77b8f5b721794903c2800b08e916757eac5e120ea840a8dfb1e0;
  assign mdsMatrix_29_8 = 255'h49d5e85b08d1240c6c43afeba84a82b43b5ad2d71238e5f1e1362d2cd27202bf;
  assign mdsMatrix_30_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_30_1 = 254'h35fbe93d76bd97506c40e9dbc3fac20c2454a3e1fd38f163a08ab68e7d1b856b;
  assign mdsMatrix_30_2 = 255'h5ef529ae0a04c4faeecb360f7533051ae7b75401c03ac5afe7bd1071fcc69646;
  assign mdsMatrix_30_3 = 255'h41522e0f2836f5012ecd0031b13cfaadd5370224b81735e41230c4210372423d;
  assign mdsMatrix_30_4 = 252'hb087e1f6c147fd2efd0dab6f95c8e4c8b937573a2dd634d962c51a1361ed41e;
  assign mdsMatrix_30_5 = 255'h43c36242c3dc4732b64b82e4bca568298f3c5ad09adc24d34aa276afe383b52a;
  assign mdsMatrix_30_6 = 255'h6cc879dac7a9cc9df41994916543897f6d5ef22e5d4ed317eabff7e0bc77dda0;
  assign mdsMatrix_30_7 = 254'h33b2b707fbbed03e6acf73ae8861e255a0b54b4c0d63fd8f690582aa3139887d;
  assign mdsMatrix_30_8 = 253'h16073337d84d3c256a405bcf452e3a1ad6004002bbd49d3ce2363a3ed1bd47cb;
  assign mdsMatrix_31_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_31_1 = 250'h340f55f485257dcc9f1bdba20dafb7b55641537dc0992e7ca67b28217aef258;
  assign mdsMatrix_31_2 = 252'hed7ab6e3a9f056345a48e26d6aef72cb36249145b8fd981d164c61a240c6e91;
  assign mdsMatrix_31_3 = 254'h3fd36f2dba03da199297f0b5b6376d4a5d8700c7925d31bd4fa8e6574029db7a;
  assign mdsMatrix_31_4 = 254'h3bc8fa13d824729b9d057bf59406fd9c9a2089e7d6830101192c39917a49137f;
  assign mdsMatrix_31_5 = 253'h1d8e67b8558d29c78e41181152a44faedb423a8754ea9ae0b90fbc761b515f54;
  assign mdsMatrix_31_6 = 255'h6205f54c7f3064ac9df7ed150f4dab4af85942be9ee8fa9c970a783704081abd;
  assign mdsMatrix_31_7 = 255'h54fa57135950320389733a7cae63890213fdd3d11845325c83e4179620f9648b;
  assign mdsMatrix_31_8 = 255'h654ae17d61d404c666a687818244eec21f49c636ec328275cca841fe2a8df05a;
  assign mdsMatrix_32_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_32_1 = 254'h20fc4af967942bd311eac60f246d2509508fcbbd13815f8c4a53e82abbc57426;
  assign mdsMatrix_32_2 = 254'h3e80f495d2a556ebe0d9177b3311cb3f36f4ea63351c88ee18137f3c34a18901;
  assign mdsMatrix_32_3 = 254'h28043951bbc4f15476f88bdd42b63be862067d138bbd3e13d6cdbc3a06ae9258;
  assign mdsMatrix_32_4 = 250'h21121b838295b025b9c0c68888b62767e1ee9b688d9062a6da427bb9cbbf801;
  assign mdsMatrix_32_5 = 255'h415ce9e487191504b37535e5ec17311239b532073feffc55a54fe6daf0b87e0e;
  assign mdsMatrix_32_6 = 254'h2d2382cf9994518bfd5646e9dd9776a63c00cb6835d8b3260688fe8a41f6587c;
  assign mdsMatrix_32_7 = 254'h3a25ac7b1d7160d13f8f997c8ebb7f6b988dbbb1393845f129eda86eeb820630;
  assign mdsMatrix_32_8 = 254'h269a43a3c86e65d7bcd8efa93906caa4c46fa4ac212aa240b5c525a9b814d9d6;
  assign mdsMatrix_33_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_33_1 = 254'h2dbe6f2067da3f73f04a6ff95a5f397b35f68808685fa12bbdb0dd0cf9ab9026;
  assign mdsMatrix_33_2 = 253'h1d919b729c6d287a18801f6ae9c6bab913b26655a5a71d6ec0e15757ed445529;
  assign mdsMatrix_33_3 = 254'h3bef316cffdf758a19c2d494acedac470f68ec245571a837d6d64891152004f3;
  assign mdsMatrix_33_4 = 255'h528ab9dc5c7e9921640e776f57db510cb358415c35b4aede1b519b3e8d1e0093;
  assign mdsMatrix_33_5 = 254'h272a81f471806b2dd05771d4ce8b3260c2d4c8a5e014b66e1c5d0314cae8046e;
  assign mdsMatrix_33_6 = 251'h4d420e6b25b5bceb08c669c228451ebef520b2a54eceec8b8eb2a791de83317;
  assign mdsMatrix_33_7 = 254'h3dcb79616a3f3b4cb2b5aa74b27d8a2cc0a7d97a626423bc625aa7a50dfe9f08;
  assign mdsMatrix_33_8 = 247'h462a7cdb5a3c1c6e67b2fabf9f4683a302938be6f432828f32064e1ec99fb5;
  assign mdsMatrix_34_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_34_1 = 255'h5ce192c585128651e2ec175e13ef0428cd477ed07cc5e3d801cf376bb7af9bad;
  assign mdsMatrix_34_2 = 255'h7275ab503c14c7e3b27b072151ccb3fd0fae9bce59bd3fe3b95bdefd99c4f5fe;
  assign mdsMatrix_34_3 = 254'h334d0a97a4d96aad5735fbab438e5757f4f92649b0de11aef748b5d3419db942;
  assign mdsMatrix_34_4 = 254'h339eb21627699a78999b0b9faf1f10ada6c6288a20ec0be5c0c730ee14a2b478;
  assign mdsMatrix_34_5 = 255'h5d13239d433b926289786f06342d6d1d953c23c22a98fb5c377267be0f5083f1;
  assign mdsMatrix_34_6 = 250'h250dec55a88d6516715ce496311ef6dc78a6175e66cdd74b9a7e58fd2aef85e;
  assign mdsMatrix_34_7 = 253'h16b1390a0af9c19f59bba840cc3edad8ffdf2eda8eddaf690052daceb5185e89;
  assign mdsMatrix_34_8 = 255'h6650657d0e89e95f9d5dc0e2929be7d5660befeb2e37808bc926601a24bb2f5f;
  assign mdsMatrix_35_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_35_1 = 252'h804bba256fe110808d100b9bdf701885604a7ce2db2ce790b48c58f43bbc3c9;
  assign mdsMatrix_35_2 = 255'h6de1d82b5299f6bb3c44b1b2a77c613bc6e6a2c9c36d99b0961c633780e7440c;
  assign mdsMatrix_35_3 = 252'h90c0fda336a7745b0807cf45b5d6d79d9f130115f610caadc786c2aaaf995e7;
  assign mdsMatrix_35_4 = 255'h6a054022c6ccd73077fb8c6c8206b49ca3f6638700b9e2dbf67b2d02d5e72c4a;
  assign mdsMatrix_35_5 = 255'h4080237b4939e82dacd03421066c6f0317256abc8de6def918fbbccb9c5565c3;
  assign mdsMatrix_35_6 = 255'h5f6e103d3a596e57fa01bb6f0790bfdb6b68b3d149997615e648e6ba2f54928b;
  assign mdsMatrix_35_7 = 252'ha3f4d2efaf617d1914a40b9457e4feb6bbd3ed08f0423afdab2a34908c88602;
  assign mdsMatrix_35_8 = 252'hb0cec59b91ab5cc2889efed977f0e32cd9b68460f3c140ea50c5e17d836b918;
  assign mdsMatrix_36_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_36_1 = 254'h221b24c784056132cc2dbaac4e014f212c8f5a66527177063854920c63f0966d;
  assign mdsMatrix_36_2 = 255'h433f656780a4c39eaa674a233aa55b05f5d51568fd8842349e9ac28211c8e50c;
  assign mdsMatrix_36_3 = 254'h2c3771de537316e719ce98648acbde764e081cf2bc24b768315c15940fc6de4e;
  assign mdsMatrix_36_4 = 254'h3352d3f61186cc2e87b53786031aea684765f707dbadb85a1520410dda1d1e28;
  assign mdsMatrix_36_5 = 254'h30196adebaf73014c28428ab4218121482382b779bb2c3739cad5549ac75025b;
  assign mdsMatrix_36_6 = 251'h5c8bf7b2f7dd1d0837cdf864bcf05d2b6f7edf32d1574bf2f228cdabc9d529c;
  assign mdsMatrix_36_7 = 253'h10e64a7a6d6c626046f0e34b7a3399803340e62ea03c301572724fa016efb228;
  assign mdsMatrix_36_8 = 253'h1f39189b0783fad0c6e6694bfb41e9adc9ca5e31d2a716eb47d601eb0cc7b7f2;
  assign mdsMatrix_37_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_37_1 = 253'h19521e10e25dac0ea8a7a5415c687f31dfa26cc0b6dcf701fa01d902e1ff3077;
  assign mdsMatrix_37_2 = 255'h5ed0ef16f406a31fad174c3b75777a539b60cd74e5f352dd34b44cddaf6fc620;
  assign mdsMatrix_37_3 = 254'h2517bf962e231da5ca1bfe161dba6c31b6bda876423bb135efb48c574cd90204;
  assign mdsMatrix_37_4 = 254'h30d30b336074f8782c09245ad06e934f4d57c21d47cb62db759ac4949ccef04e;
  assign mdsMatrix_37_5 = 254'h2b5dc2c32c7f107d52ed1f3072c7450ac153aed91056af3804ac43e5bd677ee5;
  assign mdsMatrix_37_6 = 255'h55bddc68fca07f642d87d708d3093b7686967eaf162d292e2c8f68effbd1bb7c;
  assign mdsMatrix_37_7 = 255'h42b855abe9671be97bffd652b0343f5423cf0fde2054fb6d35cbcb0193489bf7;
  assign mdsMatrix_37_8 = 255'h48733fcbd7117d447585bfdf3bde5f4f7dc84fd9f1be13523e47ee2d2e5a0b27;
  assign mdsMatrix_38_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_38_1 = 253'h17ad2c9f333d220b1a87fc197fcea13fe5e90ef63a4e909d949a72af2e81489f;
  assign mdsMatrix_38_2 = 255'h618fae4f9f0947b2cc8d4712918db0d2714d12a8e3a550a7bfa7b87df5001c3f;
  assign mdsMatrix_38_3 = 255'h4cfb214582ca64600912e52df150bba8657ae8160d2224fed1eee109069a49fc;
  assign mdsMatrix_38_4 = 255'h66eaf3ac6adcb1a86d1fe25190b3f0a4b871eb67ece466802fe3fd6a5c345f04;
  assign mdsMatrix_38_5 = 254'h296bddae2f692643e9253f3869286aa0595275ae191ccbe0d42bf352eeaa98b2;
  assign mdsMatrix_38_6 = 253'h196035b2ff805e71bf6b36b98d3ae139608c297e639ab62cc020bff04e95c217;
  assign mdsMatrix_38_7 = 250'h35e3bfa30095dbc57d630e280dde652c8bf4e53c8c13c59d5a98aef519d3ec2;
  assign mdsMatrix_38_8 = 254'h3c00d5a12f8fc3cf0b8111329f6c7ad38b64c6772cbc410fdca9b9f050924fb1;
  assign mdsMatrix_39_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_39_1 = 254'h290aff34e9317863f74cf584b33937410f1838752504cba3e24cb1c4f4643c84;
  assign mdsMatrix_39_2 = 253'h1ca4945f7f39eac7617f36578a89ecdbf49afad3ad5214a67b63d6eb22f30745;
  assign mdsMatrix_39_3 = 255'h6daa9779ad9724ce2183bfea5f6ade167c5c3f0c9b34e801ec0e1fb20d9d1d29;
  assign mdsMatrix_39_4 = 255'h72eb448211ca3c6d93763292688d8b2ca4a0e3c2ce1c0d4c8929c9f0c0e1cf2a;
  assign mdsMatrix_39_5 = 254'h35f797035427b3f6cde0d9bc2152a2ce142072a5899e8957b494612e8c32a6a6;
  assign mdsMatrix_39_6 = 252'heb4cc131a6e5815b57ab853367005cd5c91e76a74faeff21bc49ed06c13da2f;
  assign mdsMatrix_39_7 = 255'h5e67c340f44d3d2c95170d4fd112d0280bffd096d3eb6a09c60e8c59be98a330;
  assign mdsMatrix_39_8 = 254'h31cf22654ef5bd147d2c723be82f03921ab0769b50a71af598b5b91b45f80b8e;
  assign mdsMatrix_40_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_40_1 = 255'h470c7780f1d9efb8eef3839542c52e79d2ea274cd20dac322c8a0a87f9806346;
  assign mdsMatrix_40_2 = 255'h4618eb35f4fe16aed6f471782141b11d296b2d8f1b4edfa8b85cda4cc5320dde;
  assign mdsMatrix_40_3 = 253'h130ed008055340555dfd15e54e177a4e2f9e0d3b8d47b677d8be5793553b7573;
  assign mdsMatrix_40_4 = 255'h557a4bbd8176fad40cc0578f941653c8d03eeb9f28d932516131ae40cedf439e;
  assign mdsMatrix_40_5 = 254'h3912604c9686811b7e50d89cd4c3969700dc3bb409a556b14582b852c75cc952;
  assign mdsMatrix_40_6 = 255'h631aff9893cd3550e648e53a86e7798aa3f6c457c2ea461100e77eeb035a1060;
  assign mdsMatrix_40_7 = 253'h1375d0002b73b0933107cd7ec60a1525d33619af78e1ffd72533ca3e5837c12c;
  assign mdsMatrix_40_8 = 250'h3c0b74f2fd93c0c011d034247e96d71b413096a21ec5c24b11c7b51abc9ea54;
  assign mdsMatrix_41_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_41_1 = 255'h72bbf33fb95bc2d48a664e3c3c38d299a9e6faa02ece3297aa3839ff891d2f3f;
  assign mdsMatrix_41_2 = 254'h3287ff0d4b06d67e24cdd2709f880809ba3479061a4e8a47e626e4a6548012bf;
  assign mdsMatrix_41_3 = 255'h71fbd49f1bccc04a7251e5259eb49b4d5a03a30148cbe75a7a21d2aba4121de5;
  assign mdsMatrix_41_4 = 252'hc14c281d194c3b436ebb2f8bf3dd74d22d589f60da438cd2647e11c9de35c9f;
  assign mdsMatrix_41_5 = 254'h3f8c4fd654df5e85e12dd6dca134b41a7c02c9644b49911ba930052d98e8dcfb;
  assign mdsMatrix_41_6 = 255'h6f514985be61d45baa2ed671691a72f4a6b64d33517b7c633ac7f56ebf3092cb;
  assign mdsMatrix_41_7 = 252'hf37b86a03567e3b137bcb5d037795a357c3585a0f48a6e14865b11277d0525b;
  assign mdsMatrix_41_8 = 255'h5bd33b5819c6be2e4bd68aedc676033cf2d74065f0de1dfb373c1e939072dab5;
  assign mdsMatrix_42_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_42_1 = 255'h6d8381b0c193bc67e9700209a1121cbea798b3777abf3af57f0298721cd108ba;
  assign mdsMatrix_42_2 = 255'h4d07f8e896b5ee22b289406785eb82509c246b7ceb10a416d05f511e185df209;
  assign mdsMatrix_42_3 = 254'h3744a21d1ec1607301dc048ba8e8e205b2783647984f62ac1a00deb806fa2bc2;
  assign mdsMatrix_42_4 = 254'h2c164d7a0f76c06706e4c92463e343ba334f8c4da1ee705b3728aa58050f2ad7;
  assign mdsMatrix_42_5 = 255'h6461107909576c46ca2fe300449111af801d56f5b81eb5977994335a726aca89;
  assign mdsMatrix_42_6 = 254'h34f07c4269feeb34d1fa0d3830ef286ed2eba687f7c89a366c2e42ccb9281562;
  assign mdsMatrix_42_7 = 253'h1f7fbd4c6028aff0054808223ce91ec285644e07a7e9d96750475b5dbece45f9;
  assign mdsMatrix_42_8 = 254'h31dd82875bfc612732ea2410d671d2a25248ecfa9a99e26b95a055247cead623;
  assign mdsMatrix_43_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_43_1 = 255'h434fd5d417f55d62e1051517454286ffd06892b02c3bdc82d807abef21149716;
  assign mdsMatrix_43_2 = 255'h4afe622d617a4bb7e6c9542c12a4361df868a75a24784357442bae23cea36334;
  assign mdsMatrix_43_3 = 255'h4b03101a7fbfd511a1b4391bdeb9c2d121fa95cf0d1dc5d746a72c1e91e5c22d;
  assign mdsMatrix_43_4 = 255'h736ac98bf915b4730b5b08cb6e4040380eea3b0f7e3e1ff96d4397598dfc7af0;
  assign mdsMatrix_43_5 = 255'h6bde018f9b73a44e6e7308dc7220d10aa364f179509e1e85e107d99ac0c80bfc;
  assign mdsMatrix_43_6 = 252'hc0efc6a4224dd789ae1937df0ead172082c06f136ecc46bad51ea33de46c506;
  assign mdsMatrix_43_7 = 252'hb04eea3fb72e3c91807a986d206e7d0b096995db0cebacc7f6585d26748f0ca;
  assign mdsMatrix_43_8 = 252'hc36717f1aabb0a7bcf2933001db3cbd669ece7db4eb197cf34581c02e9bd476;
  assign mdsMatrix_44_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_44_1 = 255'h6dd7aaf471a7c6f77daf583495e675a6ad087b5b1e8fd495639ba381d688897a;
  assign mdsMatrix_44_2 = 254'h29f0ff1f8ec75534a7de2ab44e8108446fe11676d4f2c6994f03bc95327d1057;
  assign mdsMatrix_44_3 = 255'h73b09cccd7d74a09bfec7e9055c571a335c17b5eb0230e6d20542ebef39e7529;
  assign mdsMatrix_44_4 = 252'h8aa496ece4355d708d2e549ff43b23c008a000e2c1454671a65f15f17900bdf;
  assign mdsMatrix_44_5 = 254'h3824cca4500baadcac35c0470ed9dcecd0c69ddd248aac7285ed157d2ce54b97;
  assign mdsMatrix_44_6 = 254'h23bd72719580cbc49c210cc1676215da1ec7262605e1895a4ff1f47c286b1540;
  assign mdsMatrix_44_7 = 254'h3ffbe7b4cc5d36c11de0168c752a3428868445078456242fccddef3359eb5840;
  assign mdsMatrix_44_8 = 255'h4ebc8de39fae1b161974d2e845d4ec3eb843aef68972d2049b7fa6959fbd58e7;
  assign mdsMatrix_45_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_45_1 = 254'h2822fe27149fbfc0ec460534ae47ec0d2dedae0589ffd81f9a252aa567f91fe5;
  assign mdsMatrix_45_2 = 253'h1c280548a4580a43b6b1d4d05d8ad40a28a79fd9c824114c23c3199148e44e6f;
  assign mdsMatrix_45_3 = 254'h270f345320bacd2b1a6080525d2baee9e4af964b75357887507bf7df9e67f025;
  assign mdsMatrix_45_4 = 254'h3f9183ca49af93e97db8f1a84b40e80c039f4124d289a43f2e08e3b0a5faa9ea;
  assign mdsMatrix_45_5 = 252'hd42cb8f9f407f1bd94894f56e9d6af2a6ccddb7bdddf62e675fecbc204a9124;
  assign mdsMatrix_45_6 = 254'h2d3db4c5c22b2055cb54e066c284dbf8c8a1af3c44d70016d7802571ba28c520;
  assign mdsMatrix_45_7 = 255'h5f3ac4cddd2221419050bc2d634568e2e2124a93442d019a76465ba0be2821c7;
  assign mdsMatrix_45_8 = 255'h56a68b51b6bcf591c47ec89a7b043cb1bf9d5933a967ac7de1bb0ddbbdb54220;
  assign mdsMatrix_46_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_46_1 = 255'h494a1e731275471636031417140cd8465fcef18a140fd144b60c28ac26f60722;
  assign mdsMatrix_46_2 = 254'h236b03f729c6955e863eb0dd4ae5eaa4460ab245c274a56a776f779f237ccbb3;
  assign mdsMatrix_46_3 = 255'h41f458fdcd0101dc37bb560d7f3196e64cda5e35e3374d18d93cf3bca91064c1;
  assign mdsMatrix_46_4 = 255'h451911ad69a54bb32c85d0736bf2b0b3e9e776181dbf80cc147da001dcefdb26;
  assign mdsMatrix_46_5 = 253'h14e644f2d9fb6c7f1aa4db5c4908b6df9044251df1c4c7720071fe82b5fcaa4f;
  assign mdsMatrix_46_6 = 254'h3abf14ee6d4c389ec931a3509202c97b896a4f212c04e24cef7191ffccafbe30;
  assign mdsMatrix_46_7 = 253'h1d6125b340e4721f959408d6d179f6421ffb918dcd6483be75a9773869df45be;
  assign mdsMatrix_46_8 = 251'h56bf317b6e109ddc731dac136bb4756c63bd46090804452e46232a079c1979e;
  assign mdsMatrix_47_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_47_1 = 254'h26470dc3aa29824d86079254da14c59a7c1f8d58b7ac7684a788bdfd04aea542;
  assign mdsMatrix_47_2 = 253'h16c87159a9cee4cc54f88a3f64846a5b176e6617dc1d30ffe37e7a4c06da4211;
  assign mdsMatrix_47_3 = 255'h4c7b59f25647fd6851eb16c738e9b1c2086e3726b93b1788cca1c241ca3ffda8;
  assign mdsMatrix_47_4 = 248'hc594eaa1ac0879d15faf16ebd3bde3abe454063289e55f5e00fb5b04278481;
  assign mdsMatrix_47_5 = 252'ha4c8c310f8f31c30ac44397d90919c2bcd2afef334a56db64ad3d1a3799bd16;
  assign mdsMatrix_47_6 = 255'h4831525f714d1e5726fcaa340c68b9f9c95a33679663a72f455c194ef2e6ce1f;
  assign mdsMatrix_47_7 = 254'h3243d900a85840b999a9ccd3e2bf35fc65b82bc5e0510d079da1a7d5ed2b8cf1;
  assign mdsMatrix_47_8 = 253'h17078f34f2f1d45917494cc110612fa588beedd8c2fab1894b8421a6d1b27065;
  assign mdsMatrix_48_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_48_1 = 255'h6bdfbcb0002b78d036ef649db17074a4d3fffc6fd3b92fddbc1237791811f73e;
  assign mdsMatrix_48_2 = 255'h573cf740a76b5393359a702382ba4a90db980966a53c6bda70539af2536626c7;
  assign mdsMatrix_48_3 = 254'h2f7f845f4dfea0a313345dc732c6ab8524f001bcd5b4714dd77be40fc50d407e;
  assign mdsMatrix_48_4 = 255'h59787396483541a87c42987718facd587724f0603bf6579e3b540dbe5060bc5d;
  assign mdsMatrix_48_5 = 255'h4f4244dd8dd24964482285b1d7dbb0ce3a4687b9427984ebfa528ccb08b6f9f9;
  assign mdsMatrix_48_6 = 254'h22a726fd8f3925e435d1c28d011cfed2653ce157e4139345f11b986ceb72a4ee;
  assign mdsMatrix_48_7 = 255'h5d17c2a47c1adf1ba57c54b37e8c5ddbb3a9598f4a8c05a5eeecbb209c83aa7e;
  assign mdsMatrix_48_8 = 252'hed5a9566256766e80abe96c0d70201f4e18364fbe5fff7d34aaf9aa3c7b96cd;
  assign mdsMatrix_49_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_49_1 = 255'h72d719b408ca4fe7541a383409f94dea05d5fbcd8fb3193ff733c373f386ede0;
  assign mdsMatrix_49_2 = 253'h1d7b1859053be2b74817d4587f148e233fd0736e9fc65b7e0497df591ca2844c;
  assign mdsMatrix_49_3 = 254'h3a8ea002e1b3e9f28509989a8487e7cacbdaa54db00e7a0b78f9554d8edc2116;
  assign mdsMatrix_49_4 = 254'h2bc15419c9f224509e9c1b357fa61f460f90825f803ca6b44cb195f978d9e852;
  assign mdsMatrix_49_5 = 249'h18441fc84626b5993c6a8afa1dd7c191ef4c4a70f91bf97e47202643a2d1e30;
  assign mdsMatrix_49_6 = 252'hf72fa00ff3aa29b03932b63a70b99531eaf6a144de1c011ce32f50d805a7edd;
  assign mdsMatrix_49_7 = 255'h5c72a2634830023150dc47a8990fe3533a91fa2ecd25de238831322d9206fe4b;
  assign mdsMatrix_49_8 = 252'hda289e60c19d342e63f946f6c4d8cd189b868603b86568e81835ab3f4bab036;
  assign mdsMatrix_50_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_50_1 = 255'h584862032ae89ec10c3db90b140d1050b296eeb0428d7f5ed61158e569be8986;
  assign mdsMatrix_50_2 = 255'h47267d748e370323ef3ffb4f8c4c3e7e452302dde41b624f0f51b79fd0eaefdb;
  assign mdsMatrix_50_3 = 251'h728c83fe4df79da243a15825a6a7cc1b02003e2a860ced660ac3ce0ec70289a;
  assign mdsMatrix_50_4 = 251'h6f23b0d0196eb3061b001a10945367f22490c269dff4356972968add3561b3d;
  assign mdsMatrix_50_5 = 255'h609a91d61ab565f8b2377bcb217fdcb6d10c56a632656a6f5c2f3f91d200e445;
  assign mdsMatrix_50_6 = 255'h666b188a4a382953e8c550c826f3869f3c0b1e6c04aca616d5667c09db5abbd7;
  assign mdsMatrix_50_7 = 252'h9edf2bae7f14200ac5df814369e72c5b61ea7749597640c809587c6d1b216c5;
  assign mdsMatrix_50_8 = 253'h1c1ff94d3bfeffb3a01dd472d45cebffe787e44c9bde14e04e5b4318d0388ea6;
  assign mdsMatrix_51_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_51_1 = 254'h2ab23626a9b2dd74fee9ad313bb74fe618e00af6617cceda0b350a61f38d08f1;
  assign mdsMatrix_51_2 = 254'h370991d29f361e5eec74dc7e2ec1fffa019d5b36dce9ba8023a02a1ba237ce8b;
  assign mdsMatrix_51_3 = 255'h71a278b2b0fa1a3bacb8657521b06a0ba2795b65ef2718a6e764dd51065a8d04;
  assign mdsMatrix_51_4 = 255'h464aa80367ca6a1b0190f3ae9306dda62bc2c5f10d787439bcfd3d4d6fe116c3;
  assign mdsMatrix_51_5 = 255'h59b45ba89c9644c803d33d65955d970bf2e09835563b52dba4a3aae6ee58cda2;
  assign mdsMatrix_51_6 = 254'h334e31a8535ebfd46052a95d7750d32e6098720cc1ce2c6dc87c826ea277a285;
  assign mdsMatrix_51_7 = 250'h21546b539b3a24cc728957d42e5bbd6e46bfa7ee350ac929634406366dba83d;
  assign mdsMatrix_51_8 = 254'h39ffcccd6c3143a1110c545561580db367a9023afea15cb797eea5e34b4179ac;
  assign mdsMatrix_52_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_52_1 = 255'h68f4fd6891cfe48ab116bdf7a98214150d99be14d27339f235fb2cea8713cd66;
  assign mdsMatrix_52_2 = 252'h830f37f0b5714f0e586ee7a1fc9ff25b8bc645df69a21963a0c10331049fe37;
  assign mdsMatrix_52_3 = 253'h125cfa3ac456c4afd030e4e2c82d0da84e6a389df7fa144763a8b77e65023b74;
  assign mdsMatrix_52_4 = 254'h37de530f854619dc75937c3baef6310b5334256c6163928c5612b472613203cd;
  assign mdsMatrix_52_5 = 255'h58c36b9f6b59f8f4fde589b58bcf0d2605c9d9e99f95ca36a9574ce8606a52fc;
  assign mdsMatrix_52_6 = 254'h322499b315811b81bb5ac39d902d41c5aa860876d4e0c8f0e56cb892f71d1ccf;
  assign mdsMatrix_52_7 = 254'h32cd9df1d750b42f2397131ccd2f5513949b25f8a6d87edc42612371f4445e1d;
  assign mdsMatrix_52_8 = 255'h5941928b0fe69f53a75fe54afad7a1cc13169040bfb0d99fea52653a2998d3a7;
  assign mdsMatrix_53_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_53_1 = 251'h5fc741f8022d460598afa8ae2b6abccf4bca2e15959d82f83cf444eeb487a6c;
  assign mdsMatrix_53_2 = 255'h58b1fb3eee9c45eb1849a5ddf3d48b7c8f80623dab42c59a771fcfb2f50edbe8;
  assign mdsMatrix_53_3 = 255'h6a7be32c6a7207166ebf7955757427b01ec37636157694100acabc08545fc582;
  assign mdsMatrix_53_4 = 255'h565b3350f47046a1cc8cbb39172e9539e47ed8a10110358e15ba1feac2715793;
  assign mdsMatrix_53_5 = 255'h5fbfa6786604596bcd03d693005bfaf4fb731072946a7b256d2e74d84b77f2e8;
  assign mdsMatrix_53_6 = 255'h4a0dedf9e2f54fd8c54ccc8fa911ea9d06803e1dd661022a39fc85484cbf36d1;
  assign mdsMatrix_53_7 = 255'h5a006823c873bc748e3dea6ad52730a519e81353b015c6a2087ac8b0a3ccab3d;
  assign mdsMatrix_53_8 = 255'h4a2c077d1c50500e829c7a1e05624161298e18e14882580e4c66e6f2d15ea5c5;
  assign mdsMatrix_54_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_54_1 = 253'h19da476a1a02265b139f9885a91cc1bdaa95e34da58d0ce1f5f5a8684ab5ce41;
  assign mdsMatrix_54_2 = 255'h4390f5bd56803f8597758e254b624d8be390375dcb652bc42071d2c314115806;
  assign mdsMatrix_54_3 = 252'h81da03d874e81ee8585b13e09d14a8f035edf2f28fb8d520e581554ae890d86;
  assign mdsMatrix_54_4 = 255'h720dad058670ba93c2bd27b373bddcb203317d43bc5ea9cf4ef409698d919e56;
  assign mdsMatrix_54_5 = 255'h47b910606fb08d4dff791ccf392fb7a3d4a112f3ae76e030c36e7740096d1d3b;
  assign mdsMatrix_54_6 = 255'h6c3de1834b5b0e65c97fee80d8aabb87d671a6a31aad80da39486fc5d7869215;
  assign mdsMatrix_54_7 = 254'h2112cae26c3e7854db8fccc291f09ba32b9a117e8b09124bc2f0798b0194facd;
  assign mdsMatrix_54_8 = 254'h3e9f940cd172a1003cb40b1ab7b476c57906c3a915972abb1fdcd49450ea8cd0;
  assign mdsMatrix_55_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_55_1 = 255'h72ca702245e2a01dddd02eec5dd3dbdfe906ca3ed933ef703014b8b1cfcd9def;
  assign mdsMatrix_55_2 = 252'h802e8814ab7b08fb04be200ba2e2a3c64d9da59ff7bc5b94773eb5116f39635;
  assign mdsMatrix_55_3 = 253'h1b908c29964179566229d9c13b26136326dd3fb509a37e829e95043afe2557e7;
  assign mdsMatrix_55_4 = 255'h49d1e759735cd0b12588076265725959f0c4c473c93ec3c310c0e4c195579d88;
  assign mdsMatrix_55_5 = 255'h71e15bea13d41f00e0ee1e0ef456183d9d4d1df01f052d27aeb29a7ed7705f19;
  assign mdsMatrix_55_6 = 255'h4828d5b47bd7159d9dbe04929c96b74af368be1c0c7d77af6e4131d7e146fb15;
  assign mdsMatrix_55_7 = 253'h17fac39793e8dd8d7a4f6c9f671d35188c0c8974ba33c662de9660f803fa99b5;
  assign mdsMatrix_55_8 = 255'h5e796584458e6a7e3dff51ab4e764831f6ebe4eea260a1efd2881a2e340e3507;
  assign mdsMatrix_56_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_56_1 = 255'h73ceab31cb0d53b6a30a68a20a8735c2532f113d3365bb520000001eccccccae;
  assign mdsMatrix_56_2 = 251'h6004d4d83630ca1d2b8ab46124b477e072c5bda77c92ca1745d168586fb5930;
  assign mdsMatrix_56_3 = 253'h12a38b6ead3faa51fd56626e70e5af085956047e1b60df3ad1745f97e8ba2c0b;
  assign mdsMatrix_56_4 = 255'h4c1014683c3771b9df0074817e18cb0cfb4761a1d77ac8b48f377a0c479bc49c;
  assign mdsMatrix_56_5 = 255'h6dbca8596bbb5645c60e1f6b728a7f66d4ca5006a7f505bc27627c8113b134ba;
  assign mdsMatrix_56_6 = 254'h3eb5fd8b2eeb0fbf8f71a437cdfc6baf60884e20d48edf109d89d3bde85e8ac8;
  assign mdsMatrix_56_7 = 254'h37ee0adb2e3052bce71d2f5b8a076c265b962f18a4e62b414ec4ee64c0fc0dab;
  assign mdsMatrix_56_8 = 254'h2ed49d9cea20f0649bedb84f5e3221d5ed1fefac01af3bf5627626ffcf593232;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign tempAddrVec_5 = io_addr_regNext_5;
  assign tempAddrVec_6 = io_addr_regNext_6;
  assign tempAddrVec_7 = io_addr_regNext_7;
  assign tempAddrVec_8 = io_addr_regNext_8;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  assign io_data_5 = _zz_mdsMem_5_port0;
  assign io_data_6 = _zz_mdsMem_6_port0;
  assign io_data_7 = _zz_mdsMem_7_port0;
  assign io_data_8 = _zz_mdsMem_8_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
    io_addr_regNext_5 <= io_addr;
    io_addr_regNext_6 <= io_addr;
    io_addr_regNext_7 <= io_addr;
    io_addr_regNext_8 <= io_addr;
  end


endmodule

module MatrixConstantMem_11 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  output     [254:0]  io_data_9,
  output     [254:0]  io_data_10,
  output     [254:0]  io_data_11,
  input      [5:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  reg        [254:0]  _zz_mdsMem_5_port0;
  reg        [254:0]  _zz_mdsMem_6_port0;
  reg        [254:0]  _zz_mdsMem_7_port0;
  reg        [254:0]  _zz_mdsMem_8_port0;
  reg        [254:0]  _zz_mdsMem_9_port0;
  reg        [254:0]  _zz_mdsMem_10_port0;
  reg        [254:0]  _zz_mdsMem_11_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire                _zz_mdsMem_5_port;
  wire                _zz_io_data_5;
  wire                _zz_mdsMem_6_port;
  wire                _zz_io_data_6;
  wire                _zz_mdsMem_7_port;
  wire                _zz_io_data_7;
  wire                _zz_mdsMem_8_port;
  wire                _zz_io_data_8;
  wire                _zz_mdsMem_9_port;
  wire                _zz_io_data_9;
  wire                _zz_mdsMem_10_port;
  wire                _zz_io_data_10;
  wire                _zz_mdsMem_11_port;
  wire                _zz_io_data_11;
  wire       [254:0]  mdsMatrix_0_0;
  wire       [253:0]  mdsMatrix_0_1;
  wire       [250:0]  mdsMatrix_0_2;
  wire       [254:0]  mdsMatrix_0_3;
  wire       [254:0]  mdsMatrix_0_4;
  wire       [252:0]  mdsMatrix_0_5;
  wire       [254:0]  mdsMatrix_0_6;
  wire       [253:0]  mdsMatrix_0_7;
  wire       [253:0]  mdsMatrix_0_8;
  wire       [253:0]  mdsMatrix_0_9;
  wire       [248:0]  mdsMatrix_0_10;
  wire       [252:0]  mdsMatrix_0_11;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [252:0]  mdsMatrix_1_1;
  wire       [252:0]  mdsMatrix_1_2;
  wire       [254:0]  mdsMatrix_1_3;
  wire       [253:0]  mdsMatrix_1_4;
  wire       [252:0]  mdsMatrix_1_5;
  wire       [254:0]  mdsMatrix_1_6;
  wire       [254:0]  mdsMatrix_1_7;
  wire       [251:0]  mdsMatrix_1_8;
  wire       [252:0]  mdsMatrix_1_9;
  wire       [251:0]  mdsMatrix_1_10;
  wire       [253:0]  mdsMatrix_1_11;
  wire       [254:0]  mdsMatrix_2_0;
  wire       [253:0]  mdsMatrix_2_1;
  wire       [254:0]  mdsMatrix_2_2;
  wire       [252:0]  mdsMatrix_2_3;
  wire       [254:0]  mdsMatrix_2_4;
  wire       [252:0]  mdsMatrix_2_5;
  wire       [253:0]  mdsMatrix_2_6;
  wire       [253:0]  mdsMatrix_2_7;
  wire       [254:0]  mdsMatrix_2_8;
  wire       [253:0]  mdsMatrix_2_9;
  wire       [249:0]  mdsMatrix_2_10;
  wire       [253:0]  mdsMatrix_2_11;
  wire       [254:0]  mdsMatrix_3_0;
  wire       [251:0]  mdsMatrix_3_1;
  wire       [254:0]  mdsMatrix_3_2;
  wire       [254:0]  mdsMatrix_3_3;
  wire       [254:0]  mdsMatrix_3_4;
  wire       [252:0]  mdsMatrix_3_5;
  wire       [254:0]  mdsMatrix_3_6;
  wire       [252:0]  mdsMatrix_3_7;
  wire       [253:0]  mdsMatrix_3_8;
  wire       [252:0]  mdsMatrix_3_9;
  wire       [253:0]  mdsMatrix_3_10;
  wire       [253:0]  mdsMatrix_3_11;
  wire       [254:0]  mdsMatrix_4_0;
  wire       [254:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [252:0]  mdsMatrix_4_3;
  wire       [253:0]  mdsMatrix_4_4;
  wire       [252:0]  mdsMatrix_4_5;
  wire       [254:0]  mdsMatrix_4_6;
  wire       [254:0]  mdsMatrix_4_7;
  wire       [254:0]  mdsMatrix_4_8;
  wire       [253:0]  mdsMatrix_4_9;
  wire       [254:0]  mdsMatrix_4_10;
  wire       [254:0]  mdsMatrix_4_11;
  wire       [254:0]  mdsMatrix_5_0;
  wire       [254:0]  mdsMatrix_5_1;
  wire       [253:0]  mdsMatrix_5_2;
  wire       [252:0]  mdsMatrix_5_3;
  wire       [251:0]  mdsMatrix_5_4;
  wire       [254:0]  mdsMatrix_5_5;
  wire       [253:0]  mdsMatrix_5_6;
  wire       [254:0]  mdsMatrix_5_7;
  wire       [254:0]  mdsMatrix_5_8;
  wire       [254:0]  mdsMatrix_5_9;
  wire       [252:0]  mdsMatrix_5_10;
  wire       [254:0]  mdsMatrix_5_11;
  wire       [254:0]  mdsMatrix_6_0;
  wire       [254:0]  mdsMatrix_6_1;
  wire       [254:0]  mdsMatrix_6_2;
  wire       [253:0]  mdsMatrix_6_3;
  wire       [253:0]  mdsMatrix_6_4;
  wire       [254:0]  mdsMatrix_6_5;
  wire       [250:0]  mdsMatrix_6_6;
  wire       [253:0]  mdsMatrix_6_7;
  wire       [254:0]  mdsMatrix_6_8;
  wire       [253:0]  mdsMatrix_6_9;
  wire       [253:0]  mdsMatrix_6_10;
  wire       [253:0]  mdsMatrix_6_11;
  wire       [254:0]  mdsMatrix_7_0;
  wire       [254:0]  mdsMatrix_7_1;
  wire       [254:0]  mdsMatrix_7_2;
  wire       [253:0]  mdsMatrix_7_3;
  wire       [254:0]  mdsMatrix_7_4;
  wire       [254:0]  mdsMatrix_7_5;
  wire       [254:0]  mdsMatrix_7_6;
  wire       [254:0]  mdsMatrix_7_7;
  wire       [253:0]  mdsMatrix_7_8;
  wire       [250:0]  mdsMatrix_7_9;
  wire       [254:0]  mdsMatrix_7_10;
  wire       [254:0]  mdsMatrix_7_11;
  wire       [254:0]  mdsMatrix_8_0;
  wire       [254:0]  mdsMatrix_8_1;
  wire       [254:0]  mdsMatrix_8_2;
  wire       [254:0]  mdsMatrix_8_3;
  wire       [254:0]  mdsMatrix_8_4;
  wire       [249:0]  mdsMatrix_8_5;
  wire       [252:0]  mdsMatrix_8_6;
  wire       [254:0]  mdsMatrix_8_7;
  wire       [253:0]  mdsMatrix_8_8;
  wire       [253:0]  mdsMatrix_8_9;
  wire       [252:0]  mdsMatrix_8_10;
  wire       [252:0]  mdsMatrix_8_11;
  wire       [254:0]  mdsMatrix_9_0;
  wire       [249:0]  mdsMatrix_9_1;
  wire       [249:0]  mdsMatrix_9_2;
  wire       [253:0]  mdsMatrix_9_3;
  wire       [254:0]  mdsMatrix_9_4;
  wire       [253:0]  mdsMatrix_9_5;
  wire       [254:0]  mdsMatrix_9_6;
  wire       [253:0]  mdsMatrix_9_7;
  wire       [250:0]  mdsMatrix_9_8;
  wire       [253:0]  mdsMatrix_9_9;
  wire       [254:0]  mdsMatrix_9_10;
  wire       [254:0]  mdsMatrix_9_11;
  wire       [254:0]  mdsMatrix_10_0;
  wire       [254:0]  mdsMatrix_10_1;
  wire       [253:0]  mdsMatrix_10_2;
  wire       [254:0]  mdsMatrix_10_3;
  wire       [254:0]  mdsMatrix_10_4;
  wire       [254:0]  mdsMatrix_10_5;
  wire       [249:0]  mdsMatrix_10_6;
  wire       [254:0]  mdsMatrix_10_7;
  wire       [252:0]  mdsMatrix_10_8;
  wire       [252:0]  mdsMatrix_10_9;
  wire       [253:0]  mdsMatrix_10_10;
  wire       [250:0]  mdsMatrix_10_11;
  wire       [254:0]  mdsMatrix_11_0;
  wire       [253:0]  mdsMatrix_11_1;
  wire       [254:0]  mdsMatrix_11_2;
  wire       [250:0]  mdsMatrix_11_3;
  wire       [253:0]  mdsMatrix_11_4;
  wire       [249:0]  mdsMatrix_11_5;
  wire       [253:0]  mdsMatrix_11_6;
  wire       [253:0]  mdsMatrix_11_7;
  wire       [254:0]  mdsMatrix_11_8;
  wire       [254:0]  mdsMatrix_11_9;
  wire       [253:0]  mdsMatrix_11_10;
  wire       [244:0]  mdsMatrix_11_11;
  wire       [254:0]  mdsMatrix_12_0;
  wire       [253:0]  mdsMatrix_12_1;
  wire       [254:0]  mdsMatrix_12_2;
  wire       [254:0]  mdsMatrix_12_3;
  wire       [254:0]  mdsMatrix_12_4;
  wire       [254:0]  mdsMatrix_12_5;
  wire       [253:0]  mdsMatrix_12_6;
  wire       [253:0]  mdsMatrix_12_7;
  wire       [254:0]  mdsMatrix_12_8;
  wire       [254:0]  mdsMatrix_12_9;
  wire       [254:0]  mdsMatrix_12_10;
  wire       [254:0]  mdsMatrix_12_11;
  wire       [254:0]  mdsMatrix_13_0;
  wire       [254:0]  mdsMatrix_13_1;
  wire       [254:0]  mdsMatrix_13_2;
  wire       [254:0]  mdsMatrix_13_3;
  wire       [252:0]  mdsMatrix_13_4;
  wire       [251:0]  mdsMatrix_13_5;
  wire       [254:0]  mdsMatrix_13_6;
  wire       [254:0]  mdsMatrix_13_7;
  wire       [254:0]  mdsMatrix_13_8;
  wire       [254:0]  mdsMatrix_13_9;
  wire       [254:0]  mdsMatrix_13_10;
  wire       [254:0]  mdsMatrix_13_11;
  wire       [254:0]  mdsMatrix_14_0;
  wire       [252:0]  mdsMatrix_14_1;
  wire       [254:0]  mdsMatrix_14_2;
  wire       [254:0]  mdsMatrix_14_3;
  wire       [253:0]  mdsMatrix_14_4;
  wire       [252:0]  mdsMatrix_14_5;
  wire       [253:0]  mdsMatrix_14_6;
  wire       [249:0]  mdsMatrix_14_7;
  wire       [252:0]  mdsMatrix_14_8;
  wire       [251:0]  mdsMatrix_14_9;
  wire       [250:0]  mdsMatrix_14_10;
  wire       [252:0]  mdsMatrix_14_11;
  wire       [254:0]  mdsMatrix_15_0;
  wire       [253:0]  mdsMatrix_15_1;
  wire       [254:0]  mdsMatrix_15_2;
  wire       [252:0]  mdsMatrix_15_3;
  wire       [252:0]  mdsMatrix_15_4;
  wire       [251:0]  mdsMatrix_15_5;
  wire       [253:0]  mdsMatrix_15_6;
  wire       [253:0]  mdsMatrix_15_7;
  wire       [250:0]  mdsMatrix_15_8;
  wire       [254:0]  mdsMatrix_15_9;
  wire       [254:0]  mdsMatrix_15_10;
  wire       [252:0]  mdsMatrix_15_11;
  wire       [254:0]  mdsMatrix_16_0;
  wire       [254:0]  mdsMatrix_16_1;
  wire       [252:0]  mdsMatrix_16_2;
  wire       [254:0]  mdsMatrix_16_3;
  wire       [253:0]  mdsMatrix_16_4;
  wire       [253:0]  mdsMatrix_16_5;
  wire       [251:0]  mdsMatrix_16_6;
  wire       [253:0]  mdsMatrix_16_7;
  wire       [252:0]  mdsMatrix_16_8;
  wire       [253:0]  mdsMatrix_16_9;
  wire       [253:0]  mdsMatrix_16_10;
  wire       [253:0]  mdsMatrix_16_11;
  wire       [254:0]  mdsMatrix_17_0;
  wire       [254:0]  mdsMatrix_17_1;
  wire       [254:0]  mdsMatrix_17_2;
  wire       [253:0]  mdsMatrix_17_3;
  wire       [253:0]  mdsMatrix_17_4;
  wire       [254:0]  mdsMatrix_17_5;
  wire       [251:0]  mdsMatrix_17_6;
  wire       [253:0]  mdsMatrix_17_7;
  wire       [254:0]  mdsMatrix_17_8;
  wire       [254:0]  mdsMatrix_17_9;
  wire       [252:0]  mdsMatrix_17_10;
  wire       [254:0]  mdsMatrix_17_11;
  wire       [254:0]  mdsMatrix_18_0;
  wire       [254:0]  mdsMatrix_18_1;
  wire       [253:0]  mdsMatrix_18_2;
  wire       [254:0]  mdsMatrix_18_3;
  wire       [252:0]  mdsMatrix_18_4;
  wire       [251:0]  mdsMatrix_18_5;
  wire       [251:0]  mdsMatrix_18_6;
  wire       [254:0]  mdsMatrix_18_7;
  wire       [254:0]  mdsMatrix_18_8;
  wire       [252:0]  mdsMatrix_18_9;
  wire       [252:0]  mdsMatrix_18_10;
  wire       [253:0]  mdsMatrix_18_11;
  wire       [254:0]  mdsMatrix_19_0;
  wire       [253:0]  mdsMatrix_19_1;
  wire       [251:0]  mdsMatrix_19_2;
  wire       [253:0]  mdsMatrix_19_3;
  wire       [253:0]  mdsMatrix_19_4;
  wire       [252:0]  mdsMatrix_19_5;
  wire       [254:0]  mdsMatrix_19_6;
  wire       [254:0]  mdsMatrix_19_7;
  wire       [254:0]  mdsMatrix_19_8;
  wire       [253:0]  mdsMatrix_19_9;
  wire       [254:0]  mdsMatrix_19_10;
  wire       [251:0]  mdsMatrix_19_11;
  wire       [254:0]  mdsMatrix_20_0;
  wire       [254:0]  mdsMatrix_20_1;
  wire       [253:0]  mdsMatrix_20_2;
  wire       [253:0]  mdsMatrix_20_3;
  wire       [254:0]  mdsMatrix_20_4;
  wire       [254:0]  mdsMatrix_20_5;
  wire       [254:0]  mdsMatrix_20_6;
  wire       [254:0]  mdsMatrix_20_7;
  wire       [252:0]  mdsMatrix_20_8;
  wire       [250:0]  mdsMatrix_20_9;
  wire       [252:0]  mdsMatrix_20_10;
  wire       [253:0]  mdsMatrix_20_11;
  wire       [254:0]  mdsMatrix_21_0;
  wire       [254:0]  mdsMatrix_21_1;
  wire       [254:0]  mdsMatrix_21_2;
  wire       [254:0]  mdsMatrix_21_3;
  wire       [252:0]  mdsMatrix_21_4;
  wire       [252:0]  mdsMatrix_21_5;
  wire       [252:0]  mdsMatrix_21_6;
  wire       [253:0]  mdsMatrix_21_7;
  wire       [250:0]  mdsMatrix_21_8;
  wire       [253:0]  mdsMatrix_21_9;
  wire       [251:0]  mdsMatrix_21_10;
  wire       [254:0]  mdsMatrix_21_11;
  wire       [254:0]  mdsMatrix_22_0;
  wire       [253:0]  mdsMatrix_22_1;
  wire       [254:0]  mdsMatrix_22_2;
  wire       [254:0]  mdsMatrix_22_3;
  wire       [250:0]  mdsMatrix_22_4;
  wire       [250:0]  mdsMatrix_22_5;
  wire       [254:0]  mdsMatrix_22_6;
  wire       [254:0]  mdsMatrix_22_7;
  wire       [252:0]  mdsMatrix_22_8;
  wire       [252:0]  mdsMatrix_22_9;
  wire       [254:0]  mdsMatrix_22_10;
  wire       [254:0]  mdsMatrix_22_11;
  wire       [254:0]  mdsMatrix_23_0;
  wire       [254:0]  mdsMatrix_23_1;
  wire       [252:0]  mdsMatrix_23_2;
  wire       [253:0]  mdsMatrix_23_3;
  wire       [254:0]  mdsMatrix_23_4;
  wire       [254:0]  mdsMatrix_23_5;
  wire       [254:0]  mdsMatrix_23_6;
  wire       [254:0]  mdsMatrix_23_7;
  wire       [249:0]  mdsMatrix_23_8;
  wire       [253:0]  mdsMatrix_23_9;
  wire       [251:0]  mdsMatrix_23_10;
  wire       [254:0]  mdsMatrix_23_11;
  wire       [254:0]  mdsMatrix_24_0;
  wire       [253:0]  mdsMatrix_24_1;
  wire       [254:0]  mdsMatrix_24_2;
  wire       [254:0]  mdsMatrix_24_3;
  wire       [254:0]  mdsMatrix_24_4;
  wire       [253:0]  mdsMatrix_24_5;
  wire       [254:0]  mdsMatrix_24_6;
  wire       [254:0]  mdsMatrix_24_7;
  wire       [254:0]  mdsMatrix_24_8;
  wire       [254:0]  mdsMatrix_24_9;
  wire       [254:0]  mdsMatrix_24_10;
  wire       [253:0]  mdsMatrix_24_11;
  wire       [254:0]  mdsMatrix_25_0;
  wire       [253:0]  mdsMatrix_25_1;
  wire       [254:0]  mdsMatrix_25_2;
  wire       [254:0]  mdsMatrix_25_3;
  wire       [254:0]  mdsMatrix_25_4;
  wire       [253:0]  mdsMatrix_25_5;
  wire       [253:0]  mdsMatrix_25_6;
  wire       [250:0]  mdsMatrix_25_7;
  wire       [254:0]  mdsMatrix_25_8;
  wire       [254:0]  mdsMatrix_25_9;
  wire       [254:0]  mdsMatrix_25_10;
  wire       [253:0]  mdsMatrix_25_11;
  wire       [254:0]  mdsMatrix_26_0;
  wire       [254:0]  mdsMatrix_26_1;
  wire       [254:0]  mdsMatrix_26_2;
  wire       [253:0]  mdsMatrix_26_3;
  wire       [253:0]  mdsMatrix_26_4;
  wire       [249:0]  mdsMatrix_26_5;
  wire       [245:0]  mdsMatrix_26_6;
  wire       [254:0]  mdsMatrix_26_7;
  wire       [254:0]  mdsMatrix_26_8;
  wire       [254:0]  mdsMatrix_26_9;
  wire       [254:0]  mdsMatrix_26_10;
  wire       [253:0]  mdsMatrix_26_11;
  wire       [254:0]  mdsMatrix_27_0;
  wire       [254:0]  mdsMatrix_27_1;
  wire       [253:0]  mdsMatrix_27_2;
  wire       [254:0]  mdsMatrix_27_3;
  wire       [253:0]  mdsMatrix_27_4;
  wire       [254:0]  mdsMatrix_27_5;
  wire       [253:0]  mdsMatrix_27_6;
  wire       [251:0]  mdsMatrix_27_7;
  wire       [252:0]  mdsMatrix_27_8;
  wire       [253:0]  mdsMatrix_27_9;
  wire       [253:0]  mdsMatrix_27_10;
  wire       [254:0]  mdsMatrix_27_11;
  wire       [254:0]  mdsMatrix_28_0;
  wire       [251:0]  mdsMatrix_28_1;
  wire       [253:0]  mdsMatrix_28_2;
  wire       [254:0]  mdsMatrix_28_3;
  wire       [252:0]  mdsMatrix_28_4;
  wire       [253:0]  mdsMatrix_28_5;
  wire       [254:0]  mdsMatrix_28_6;
  wire       [253:0]  mdsMatrix_28_7;
  wire       [252:0]  mdsMatrix_28_8;
  wire       [254:0]  mdsMatrix_28_9;
  wire       [254:0]  mdsMatrix_28_10;
  wire       [247:0]  mdsMatrix_28_11;
  wire       [254:0]  mdsMatrix_29_0;
  wire       [251:0]  mdsMatrix_29_1;
  wire       [253:0]  mdsMatrix_29_2;
  wire       [254:0]  mdsMatrix_29_3;
  wire       [254:0]  mdsMatrix_29_4;
  wire       [254:0]  mdsMatrix_29_5;
  wire       [253:0]  mdsMatrix_29_6;
  wire       [254:0]  mdsMatrix_29_7;
  wire       [252:0]  mdsMatrix_29_8;
  wire       [254:0]  mdsMatrix_29_9;
  wire       [253:0]  mdsMatrix_29_10;
  wire       [252:0]  mdsMatrix_29_11;
  wire       [254:0]  mdsMatrix_30_0;
  wire       [254:0]  mdsMatrix_30_1;
  wire       [253:0]  mdsMatrix_30_2;
  wire       [254:0]  mdsMatrix_30_3;
  wire       [253:0]  mdsMatrix_30_4;
  wire       [252:0]  mdsMatrix_30_5;
  wire       [251:0]  mdsMatrix_30_6;
  wire       [248:0]  mdsMatrix_30_7;
  wire       [254:0]  mdsMatrix_30_8;
  wire       [252:0]  mdsMatrix_30_9;
  wire       [254:0]  mdsMatrix_30_10;
  wire       [252:0]  mdsMatrix_30_11;
  wire       [254:0]  mdsMatrix_31_0;
  wire       [252:0]  mdsMatrix_31_1;
  wire       [254:0]  mdsMatrix_31_2;
  wire       [254:0]  mdsMatrix_31_3;
  wire       [254:0]  mdsMatrix_31_4;
  wire       [250:0]  mdsMatrix_31_5;
  wire       [252:0]  mdsMatrix_31_6;
  wire       [253:0]  mdsMatrix_31_7;
  wire       [253:0]  mdsMatrix_31_8;
  wire       [253:0]  mdsMatrix_31_9;
  wire       [254:0]  mdsMatrix_31_10;
  wire       [254:0]  mdsMatrix_31_11;
  wire       [254:0]  mdsMatrix_32_0;
  wire       [254:0]  mdsMatrix_32_1;
  wire       [253:0]  mdsMatrix_32_2;
  wire       [254:0]  mdsMatrix_32_3;
  wire       [253:0]  mdsMatrix_32_4;
  wire       [253:0]  mdsMatrix_32_5;
  wire       [251:0]  mdsMatrix_32_6;
  wire       [253:0]  mdsMatrix_32_7;
  wire       [253:0]  mdsMatrix_32_8;
  wire       [252:0]  mdsMatrix_32_9;
  wire       [253:0]  mdsMatrix_32_10;
  wire       [253:0]  mdsMatrix_32_11;
  wire       [254:0]  mdsMatrix_33_0;
  wire       [252:0]  mdsMatrix_33_1;
  wire       [254:0]  mdsMatrix_33_2;
  wire       [254:0]  mdsMatrix_33_3;
  wire       [253:0]  mdsMatrix_33_4;
  wire       [254:0]  mdsMatrix_33_5;
  wire       [251:0]  mdsMatrix_33_6;
  wire       [252:0]  mdsMatrix_33_7;
  wire       [254:0]  mdsMatrix_33_8;
  wire       [253:0]  mdsMatrix_33_9;
  wire       [253:0]  mdsMatrix_33_10;
  wire       [254:0]  mdsMatrix_33_11;
  wire       [254:0]  mdsMatrix_34_0;
  wire       [253:0]  mdsMatrix_34_1;
  wire       [254:0]  mdsMatrix_34_2;
  wire       [250:0]  mdsMatrix_34_3;
  wire       [254:0]  mdsMatrix_34_4;
  wire       [254:0]  mdsMatrix_34_5;
  wire       [252:0]  mdsMatrix_34_6;
  wire       [254:0]  mdsMatrix_34_7;
  wire       [249:0]  mdsMatrix_34_8;
  wire       [254:0]  mdsMatrix_34_9;
  wire       [253:0]  mdsMatrix_34_10;
  wire       [254:0]  mdsMatrix_34_11;
  wire       [254:0]  mdsMatrix_35_0;
  wire       [254:0]  mdsMatrix_35_1;
  wire       [252:0]  mdsMatrix_35_2;
  wire       [253:0]  mdsMatrix_35_3;
  wire       [254:0]  mdsMatrix_35_4;
  wire       [253:0]  mdsMatrix_35_5;
  wire       [250:0]  mdsMatrix_35_6;
  wire       [252:0]  mdsMatrix_35_7;
  wire       [250:0]  mdsMatrix_35_8;
  wire       [253:0]  mdsMatrix_35_9;
  wire       [251:0]  mdsMatrix_35_10;
  wire       [251:0]  mdsMatrix_35_11;
  wire       [254:0]  mdsMatrix_36_0;
  wire       [254:0]  mdsMatrix_36_1;
  wire       [251:0]  mdsMatrix_36_2;
  wire       [254:0]  mdsMatrix_36_3;
  wire       [254:0]  mdsMatrix_36_4;
  wire       [251:0]  mdsMatrix_36_5;
  wire       [253:0]  mdsMatrix_36_6;
  wire       [252:0]  mdsMatrix_36_7;
  wire       [252:0]  mdsMatrix_36_8;
  wire       [254:0]  mdsMatrix_36_9;
  wire       [254:0]  mdsMatrix_36_10;
  wire       [253:0]  mdsMatrix_36_11;
  wire       [254:0]  mdsMatrix_37_0;
  wire       [253:0]  mdsMatrix_37_1;
  wire       [254:0]  mdsMatrix_37_2;
  wire       [254:0]  mdsMatrix_37_3;
  wire       [253:0]  mdsMatrix_37_4;
  wire       [252:0]  mdsMatrix_37_5;
  wire       [251:0]  mdsMatrix_37_6;
  wire       [254:0]  mdsMatrix_37_7;
  wire       [254:0]  mdsMatrix_37_8;
  wire       [254:0]  mdsMatrix_37_9;
  wire       [249:0]  mdsMatrix_37_10;
  wire       [250:0]  mdsMatrix_37_11;
  wire       [254:0]  mdsMatrix_38_0;
  wire       [254:0]  mdsMatrix_38_1;
  wire       [254:0]  mdsMatrix_38_2;
  wire       [253:0]  mdsMatrix_38_3;
  wire       [254:0]  mdsMatrix_38_4;
  wire       [253:0]  mdsMatrix_38_5;
  wire       [252:0]  mdsMatrix_38_6;
  wire       [254:0]  mdsMatrix_38_7;
  wire       [253:0]  mdsMatrix_38_8;
  wire       [254:0]  mdsMatrix_38_9;
  wire       [254:0]  mdsMatrix_38_10;
  wire       [253:0]  mdsMatrix_38_11;
  wire       [254:0]  mdsMatrix_39_0;
  wire       [254:0]  mdsMatrix_39_1;
  wire       [253:0]  mdsMatrix_39_2;
  wire       [251:0]  mdsMatrix_39_3;
  wire       [251:0]  mdsMatrix_39_4;
  wire       [254:0]  mdsMatrix_39_5;
  wire       [254:0]  mdsMatrix_39_6;
  wire       [254:0]  mdsMatrix_39_7;
  wire       [248:0]  mdsMatrix_39_8;
  wire       [253:0]  mdsMatrix_39_9;
  wire       [251:0]  mdsMatrix_39_10;
  wire       [246:0]  mdsMatrix_39_11;
  wire       [254:0]  mdsMatrix_40_0;
  wire       [254:0]  mdsMatrix_40_1;
  wire       [253:0]  mdsMatrix_40_2;
  wire       [253:0]  mdsMatrix_40_3;
  wire       [252:0]  mdsMatrix_40_4;
  wire       [251:0]  mdsMatrix_40_5;
  wire       [251:0]  mdsMatrix_40_6;
  wire       [253:0]  mdsMatrix_40_7;
  wire       [252:0]  mdsMatrix_40_8;
  wire       [252:0]  mdsMatrix_40_9;
  wire       [254:0]  mdsMatrix_40_10;
  wire       [252:0]  mdsMatrix_40_11;
  wire       [254:0]  mdsMatrix_41_0;
  wire       [253:0]  mdsMatrix_41_1;
  wire       [254:0]  mdsMatrix_41_2;
  wire       [254:0]  mdsMatrix_41_3;
  wire       [253:0]  mdsMatrix_41_4;
  wire       [253:0]  mdsMatrix_41_5;
  wire       [254:0]  mdsMatrix_41_6;
  wire       [253:0]  mdsMatrix_41_7;
  wire       [254:0]  mdsMatrix_41_8;
  wire       [252:0]  mdsMatrix_41_9;
  wire       [254:0]  mdsMatrix_41_10;
  wire       [254:0]  mdsMatrix_41_11;
  wire       [254:0]  mdsMatrix_42_0;
  wire       [253:0]  mdsMatrix_42_1;
  wire       [253:0]  mdsMatrix_42_2;
  wire       [252:0]  mdsMatrix_42_3;
  wire       [254:0]  mdsMatrix_42_4;
  wire       [254:0]  mdsMatrix_42_5;
  wire       [250:0]  mdsMatrix_42_6;
  wire       [254:0]  mdsMatrix_42_7;
  wire       [253:0]  mdsMatrix_42_8;
  wire       [254:0]  mdsMatrix_42_9;
  wire       [252:0]  mdsMatrix_42_10;
  wire       [254:0]  mdsMatrix_42_11;
  wire       [254:0]  mdsMatrix_43_0;
  wire       [254:0]  mdsMatrix_43_1;
  wire       [254:0]  mdsMatrix_43_2;
  wire       [254:0]  mdsMatrix_43_3;
  wire       [254:0]  mdsMatrix_43_4;
  wire       [254:0]  mdsMatrix_43_5;
  wire       [249:0]  mdsMatrix_43_6;
  wire       [254:0]  mdsMatrix_43_7;
  wire       [253:0]  mdsMatrix_43_8;
  wire       [248:0]  mdsMatrix_43_9;
  wire       [254:0]  mdsMatrix_43_10;
  wire       [253:0]  mdsMatrix_43_11;
  wire       [254:0]  mdsMatrix_44_0;
  wire       [252:0]  mdsMatrix_44_1;
  wire       [253:0]  mdsMatrix_44_2;
  wire       [254:0]  mdsMatrix_44_3;
  wire       [253:0]  mdsMatrix_44_4;
  wire       [254:0]  mdsMatrix_44_5;
  wire       [252:0]  mdsMatrix_44_6;
  wire       [254:0]  mdsMatrix_44_7;
  wire       [251:0]  mdsMatrix_44_8;
  wire       [253:0]  mdsMatrix_44_9;
  wire       [251:0]  mdsMatrix_44_10;
  wire       [254:0]  mdsMatrix_44_11;
  wire       [254:0]  mdsMatrix_45_0;
  wire       [252:0]  mdsMatrix_45_1;
  wire       [252:0]  mdsMatrix_45_2;
  wire       [254:0]  mdsMatrix_45_3;
  wire       [252:0]  mdsMatrix_45_4;
  wire       [250:0]  mdsMatrix_45_5;
  wire       [254:0]  mdsMatrix_45_6;
  wire       [253:0]  mdsMatrix_45_7;
  wire       [254:0]  mdsMatrix_45_8;
  wire       [252:0]  mdsMatrix_45_9;
  wire       [254:0]  mdsMatrix_45_10;
  wire       [254:0]  mdsMatrix_45_11;
  wire       [254:0]  mdsMatrix_46_0;
  wire       [251:0]  mdsMatrix_46_1;
  wire       [254:0]  mdsMatrix_46_2;
  wire       [253:0]  mdsMatrix_46_3;
  wire       [254:0]  mdsMatrix_46_4;
  wire       [254:0]  mdsMatrix_46_5;
  wire       [252:0]  mdsMatrix_46_6;
  wire       [252:0]  mdsMatrix_46_7;
  wire       [252:0]  mdsMatrix_46_8;
  wire       [254:0]  mdsMatrix_46_9;
  wire       [254:0]  mdsMatrix_46_10;
  wire       [254:0]  mdsMatrix_46_11;
  wire       [254:0]  mdsMatrix_47_0;
  wire       [253:0]  mdsMatrix_47_1;
  wire       [252:0]  mdsMatrix_47_2;
  wire       [254:0]  mdsMatrix_47_3;
  wire       [254:0]  mdsMatrix_47_4;
  wire       [253:0]  mdsMatrix_47_5;
  wire       [252:0]  mdsMatrix_47_6;
  wire       [254:0]  mdsMatrix_47_7;
  wire       [254:0]  mdsMatrix_47_8;
  wire       [248:0]  mdsMatrix_47_9;
  wire       [254:0]  mdsMatrix_47_10;
  wire       [254:0]  mdsMatrix_47_11;
  wire       [254:0]  mdsMatrix_48_0;
  wire       [254:0]  mdsMatrix_48_1;
  wire       [254:0]  mdsMatrix_48_2;
  wire       [252:0]  mdsMatrix_48_3;
  wire       [254:0]  mdsMatrix_48_4;
  wire       [254:0]  mdsMatrix_48_5;
  wire       [251:0]  mdsMatrix_48_6;
  wire       [254:0]  mdsMatrix_48_7;
  wire       [254:0]  mdsMatrix_48_8;
  wire       [254:0]  mdsMatrix_48_9;
  wire       [254:0]  mdsMatrix_48_10;
  wire       [254:0]  mdsMatrix_48_11;
  wire       [254:0]  mdsMatrix_49_0;
  wire       [250:0]  mdsMatrix_49_1;
  wire       [254:0]  mdsMatrix_49_2;
  wire       [254:0]  mdsMatrix_49_3;
  wire       [254:0]  mdsMatrix_49_4;
  wire       [253:0]  mdsMatrix_49_5;
  wire       [254:0]  mdsMatrix_49_6;
  wire       [250:0]  mdsMatrix_49_7;
  wire       [253:0]  mdsMatrix_49_8;
  wire       [254:0]  mdsMatrix_49_9;
  wire       [251:0]  mdsMatrix_49_10;
  wire       [254:0]  mdsMatrix_49_11;
  wire       [254:0]  mdsMatrix_50_0;
  wire       [254:0]  mdsMatrix_50_1;
  wire       [253:0]  mdsMatrix_50_2;
  wire       [254:0]  mdsMatrix_50_3;
  wire       [254:0]  mdsMatrix_50_4;
  wire       [251:0]  mdsMatrix_50_5;
  wire       [254:0]  mdsMatrix_50_6;
  wire       [254:0]  mdsMatrix_50_7;
  wire       [252:0]  mdsMatrix_50_8;
  wire       [252:0]  mdsMatrix_50_9;
  wire       [254:0]  mdsMatrix_50_10;
  wire       [254:0]  mdsMatrix_50_11;
  wire       [254:0]  mdsMatrix_51_0;
  wire       [254:0]  mdsMatrix_51_1;
  wire       [254:0]  mdsMatrix_51_2;
  wire       [253:0]  mdsMatrix_51_3;
  wire       [254:0]  mdsMatrix_51_4;
  wire       [252:0]  mdsMatrix_51_5;
  wire       [254:0]  mdsMatrix_51_6;
  wire       [254:0]  mdsMatrix_51_7;
  wire       [253:0]  mdsMatrix_51_8;
  wire       [254:0]  mdsMatrix_51_9;
  wire       [253:0]  mdsMatrix_51_10;
  wire       [254:0]  mdsMatrix_51_11;
  wire       [254:0]  mdsMatrix_52_0;
  wire       [254:0]  mdsMatrix_52_1;
  wire       [253:0]  mdsMatrix_52_2;
  wire       [253:0]  mdsMatrix_52_3;
  wire       [252:0]  mdsMatrix_52_4;
  wire       [253:0]  mdsMatrix_52_5;
  wire       [254:0]  mdsMatrix_52_6;
  wire       [254:0]  mdsMatrix_52_7;
  wire       [253:0]  mdsMatrix_52_8;
  wire       [254:0]  mdsMatrix_52_9;
  wire       [243:0]  mdsMatrix_52_10;
  wire       [254:0]  mdsMatrix_52_11;
  wire       [254:0]  mdsMatrix_53_0;
  wire       [254:0]  mdsMatrix_53_1;
  wire       [252:0]  mdsMatrix_53_2;
  wire       [254:0]  mdsMatrix_53_3;
  wire       [250:0]  mdsMatrix_53_4;
  wire       [253:0]  mdsMatrix_53_5;
  wire       [253:0]  mdsMatrix_53_6;
  wire       [248:0]  mdsMatrix_53_7;
  wire       [252:0]  mdsMatrix_53_8;
  wire       [251:0]  mdsMatrix_53_9;
  wire       [254:0]  mdsMatrix_53_10;
  wire       [254:0]  mdsMatrix_53_11;
  wire       [254:0]  mdsMatrix_54_0;
  wire       [253:0]  mdsMatrix_54_1;
  wire       [254:0]  mdsMatrix_54_2;
  wire       [253:0]  mdsMatrix_54_3;
  wire       [251:0]  mdsMatrix_54_4;
  wire       [253:0]  mdsMatrix_54_5;
  wire       [253:0]  mdsMatrix_54_6;
  wire       [254:0]  mdsMatrix_54_7;
  wire       [254:0]  mdsMatrix_54_8;
  wire       [252:0]  mdsMatrix_54_9;
  wire       [254:0]  mdsMatrix_54_10;
  wire       [253:0]  mdsMatrix_54_11;
  wire       [254:0]  mdsMatrix_55_0;
  wire       [253:0]  mdsMatrix_55_1;
  wire       [254:0]  mdsMatrix_55_2;
  wire       [253:0]  mdsMatrix_55_3;
  wire       [254:0]  mdsMatrix_55_4;
  wire       [254:0]  mdsMatrix_55_5;
  wire       [253:0]  mdsMatrix_55_6;
  wire       [253:0]  mdsMatrix_55_7;
  wire       [253:0]  mdsMatrix_55_8;
  wire       [251:0]  mdsMatrix_55_9;
  wire       [254:0]  mdsMatrix_55_10;
  wire       [254:0]  mdsMatrix_55_11;
  wire       [254:0]  mdsMatrix_56_0;
  wire       [254:0]  mdsMatrix_56_1;
  wire       [253:0]  mdsMatrix_56_2;
  wire       [254:0]  mdsMatrix_56_3;
  wire       [252:0]  mdsMatrix_56_4;
  wire       [253:0]  mdsMatrix_56_5;
  wire       [254:0]  mdsMatrix_56_6;
  wire       [252:0]  mdsMatrix_56_7;
  wire       [253:0]  mdsMatrix_56_8;
  wire       [254:0]  mdsMatrix_56_9;
  wire       [252:0]  mdsMatrix_56_10;
  wire       [250:0]  mdsMatrix_56_11;
  wire       [5:0]    tempAddrVec_0;
  wire       [5:0]    tempAddrVec_1;
  wire       [5:0]    tempAddrVec_2;
  wire       [5:0]    tempAddrVec_3;
  wire       [5:0]    tempAddrVec_4;
  wire       [5:0]    tempAddrVec_5;
  wire       [5:0]    tempAddrVec_6;
  wire       [5:0]    tempAddrVec_7;
  wire       [5:0]    tempAddrVec_8;
  wire       [5:0]    tempAddrVec_9;
  wire       [5:0]    tempAddrVec_10;
  wire       [5:0]    tempAddrVec_11;
  reg        [5:0]    io_addr_regNext;
  reg        [5:0]    io_addr_regNext_1;
  reg        [5:0]    io_addr_regNext_2;
  reg        [5:0]    io_addr_regNext_3;
  reg        [5:0]    io_addr_regNext_4;
  reg        [5:0]    io_addr_regNext_5;
  reg        [5:0]    io_addr_regNext_6;
  reg        [5:0]    io_addr_regNext_7;
  reg        [5:0]    io_addr_regNext_8;
  reg        [5:0]    io_addr_regNext_9;
  reg        [5:0]    io_addr_regNext_10;
  reg        [5:0]    io_addr_regNext_11;
  reg [254:0] mdsMem_0 [0:56];
  reg [254:0] mdsMem_1 [0:56];
  reg [254:0] mdsMem_2 [0:56];
  reg [254:0] mdsMem_3 [0:56];
  reg [254:0] mdsMem_4 [0:56];
  reg [254:0] mdsMem_5 [0:56];
  reg [254:0] mdsMem_6 [0:56];
  reg [254:0] mdsMem_7 [0:56];
  reg [254:0] mdsMem_8 [0:56];
  reg [254:0] mdsMem_9 [0:56];
  reg [254:0] mdsMem_10 [0:56];
  reg [254:0] mdsMem_11 [0:56];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  assign _zz_io_data_5 = 1'b1;
  assign _zz_io_data_6 = 1'b1;
  assign _zz_io_data_7 = 1'b1;
  assign _zz_io_data_8 = 1'b1;
  assign _zz_io_data_9 = 1'b1;
  assign _zz_io_data_10 = 1'b1;
  assign _zz_io_data_11 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_5.bin",mdsMem_5);
  end
  always @(posedge clk) begin
    if(_zz_io_data_5) begin
      _zz_mdsMem_5_port0 <= mdsMem_5[tempAddrVec_5];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_6.bin",mdsMem_6);
  end
  always @(posedge clk) begin
    if(_zz_io_data_6) begin
      _zz_mdsMem_6_port0 <= mdsMem_6[tempAddrVec_6];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_7.bin",mdsMem_7);
  end
  always @(posedge clk) begin
    if(_zz_io_data_7) begin
      _zz_mdsMem_7_port0 <= mdsMem_7[tempAddrVec_7];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_8.bin",mdsMem_8);
  end
  always @(posedge clk) begin
    if(_zz_io_data_8) begin
      _zz_mdsMem_8_port0 <= mdsMem_8[tempAddrVec_8];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_9.bin",mdsMem_9);
  end
  always @(posedge clk) begin
    if(_zz_io_data_9) begin
      _zz_mdsMem_9_port0 <= mdsMem_9[tempAddrVec_9];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_10.bin",mdsMem_10);
  end
  always @(posedge clk) begin
    if(_zz_io_data_10) begin
      _zz_mdsMem_10_port0 <= mdsMem_10[tempAddrVec_10];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_25_mdsMem_11.bin",mdsMem_11);
  end
  always @(posedge clk) begin
    if(_zz_io_data_11) begin
      _zz_mdsMem_11_port0 <= mdsMem_11[tempAddrVec_11];
    end
  end

  assign mdsMatrix_0_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_0_1 = 254'h302c90931849efc2063c4eea88a6f28e255ccc4c0296832db3c174770e25ebae;
  assign mdsMatrix_0_2 = 251'h6b410ec5952b5f1514a562da981c03f90989311ddef75e0e8e85188da845b23;
  assign mdsMatrix_0_3 = 255'h4481ea187d82cd5dfbe7dc3e7d8577db59f131249008a448ef899f34dd1e777a;
  assign mdsMatrix_0_4 = 255'h59f8cc5fbabb65875fa91aaf0fcde1d84ebdd3512912fd64b5942d4c89de12e9;
  assign mdsMatrix_0_5 = 253'h1227611d582b0856d6ec61d1aa8dfdf383f67f67c974c92dbbcdcaacab75512b;
  assign mdsMatrix_0_6 = 255'h5b65a38bba37d3a1330f0cf512779f71e4d52760a886d754a34aafb465aa8475;
  assign mdsMatrix_0_7 = 254'h34f04936ea303ee53298f304a9e3cdef1e707a57b402bea622eda672bc1d3824;
  assign mdsMatrix_0_8 = 254'h3a70206660b363944bbff71d8e2f60b5833839b0972578e372a4ff21acb15389;
  assign mdsMatrix_0_9 = 254'h271021d40a1df436a7e3e8011b0e9eda1ff53ba26714beeba3dbf8ff7e9d2709;
  assign mdsMatrix_0_10 = 249'h1c74c9ac4e56db7a1ba3e1f88535aec90990c778d538dbf4c164ee9c7309601;
  assign mdsMatrix_0_11 = 253'h158872db2fad1e085d5f479aaa41645495350a30a3bcf81db2ae283b32a66a8f;
  assign mdsMatrix_1_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_1_1 = 253'h148baf54667ffed7d4d90d898b9e977d302bd27b78c502c39397718d2197c6e9;
  assign mdsMatrix_1_2 = 253'h14d02abdfdf4c3dce8526516f2f90a7370eed2e9bf55d222843ef60487e3812d;
  assign mdsMatrix_1_3 = 255'h4ffa16c69d944a4dd61aec539cadd03574c6e9797769c8702db80284a00cc6c1;
  assign mdsMatrix_1_4 = 254'h3c8298bac6f71b1a9c5dd9f87ed63d1ea42c3bd99331ba7533a715bb8aa00344;
  assign mdsMatrix_1_5 = 253'h170c2174f6066552ed1521aca358977ecb12c508ed4c542846d5fcddd3b58105;
  assign mdsMatrix_1_6 = 255'h6b432af1c1ce6acec011809253e33da03f9a236449c754c6cd9d36d160fef9a8;
  assign mdsMatrix_1_7 = 255'h4424d7aea9cfb6b2b09db7b93fc19f56ea2dce3c04192949f4c2d520eb3eaeec;
  assign mdsMatrix_1_8 = 252'hbf9b12e0c594701454477b4042ffdf6724d62244267c19b37c61287b5556ecf;
  assign mdsMatrix_1_9 = 253'h1cab0792281bcff89a00eb5cae776b4d8ccba96d78e150ae9dc5b2620a544d9a;
  assign mdsMatrix_1_10 = 252'he29c75407df9f4211ca95238d377997a669445ccb73bbfddeea8432fae5c0c2;
  assign mdsMatrix_1_11 = 254'h2dd16090328fd6c516ed3b4208cef43624d29c89f7f74f2d2bb92920b23b258e;
  assign mdsMatrix_2_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_2_1 = 254'h29b6e416e2ca06df7b354a1b46eefbe94c1a21e8620ca65098c8d3fb3513dff3;
  assign mdsMatrix_2_2 = 255'h684090e1f5f781771efb3d640236389c699795ac4619bab832f5f24d5cc2d144;
  assign mdsMatrix_2_3 = 253'h14e5168a100c3f68a702d48510ba2315b7145225051abd421a6e8ca336331e77;
  assign mdsMatrix_2_4 = 255'h607678299dfa2751fce8684309c34873cb80122bffa214ab7885b05911b50088;
  assign mdsMatrix_2_5 = 253'h1458a110fce5c0f9557ee78ee88277f1e824fa1eef214d43014aa4e70532b028;
  assign mdsMatrix_2_6 = 254'h22e0ef8d2a55dd52e10d0701d697a5a488eae1ebf703b81cbdef74903213a83c;
  assign mdsMatrix_2_7 = 254'h2dbc1fb702ee495f04340d491bcaff9e89033958457aa7202e318d476855c9b7;
  assign mdsMatrix_2_8 = 255'h409ba307693de1af0e4f52ddd4e661f3dde3f44ee675156e33fa20556a1e8ea3;
  assign mdsMatrix_2_9 = 254'h2d511a9f07fda230e4c9ae262c56fc761b8f10099f36ea0e8e9cff6675c5f6ed;
  assign mdsMatrix_2_10 = 250'h396853561106196a105a19ec339a7f3393c46ea5af73da22cfc3205bb9c7e44;
  assign mdsMatrix_2_11 = 254'h34cdd2d620d22edcc43addf369166e31013868cab60eca08d55717106c6b97a5;
  assign mdsMatrix_3_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_3_1 = 252'hfcf50fdb0e589c51f71db6dd5b091424f7fe2ab3e6a8ad1feadd8030be10b8d;
  assign mdsMatrix_3_2 = 255'h4654bc40ef6fa78233811db264e99af771193c375cde88e42fb5b4dd6016511d;
  assign mdsMatrix_3_3 = 255'h6a3b0bd04558e97886c1144a9cdddc58551bc4fb6906c9a97cf1be01819bd84f;
  assign mdsMatrix_3_4 = 255'h5a7d2fbc5aa09233fed3a33f19fb96e463b4e10c90cd996cd0c2b6ca7a47b0c5;
  assign mdsMatrix_3_5 = 253'h1d833da2a553c5a44f6705de296f1c422fbfd3e4353945cdab6e63479f8bf8a4;
  assign mdsMatrix_3_6 = 255'h5cd2c382955beb0fd150628d1ab88407d46190ff4aaab4fb1fc29e53c13f8f3c;
  assign mdsMatrix_3_7 = 253'h1c9e96722a82c69188c071d3050b7afff1d18da665028c1b1980f46ce1ddcd2a;
  assign mdsMatrix_3_8 = 254'h30491c4ff3c5047b60b75bc14d4086b1b5eb26b41ed1df923bf05a0b42df477e;
  assign mdsMatrix_3_9 = 253'h144ea74380ef7189ab8466873bc7670da0103f22b2a09a9bb56d605bc9420276;
  assign mdsMatrix_3_10 = 254'h3450ee4b37f078f40885ba2ae4ab4061694a00054068fefca602a2bfd18304be;
  assign mdsMatrix_3_11 = 254'h2e805367685a4a0288b871067751c24b5c71389a658d6e78b3effaab37227556;
  assign mdsMatrix_4_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_4_1 = 255'h61401ccbee9e310225dd57865bbae806dc0083c042350ef205c19bd17353a759;
  assign mdsMatrix_4_2 = 255'h430098c55bdd4bdcbfe5ea4b8f9890adaf8936528e91f5fb5541603781f7c6a3;
  assign mdsMatrix_4_3 = 253'h1326d98b44fc2d75cc22e91fd1dd6a525b4aa35cb238d04f663406b72c8892d3;
  assign mdsMatrix_4_4 = 254'h38e82ff1ded664c731ef9ba33e7a8114229847b05fb8a99c4c320c477da5cb5b;
  assign mdsMatrix_4_5 = 253'h1c5f713677b5bd70e67ad3293a06b65885712cee0c4789cc1fece45f084f4451;
  assign mdsMatrix_4_6 = 255'h5c1351a24855868b8b0d82921ccc7f43d03a11d05647c5a4baaddfc02281079b;
  assign mdsMatrix_4_7 = 255'h46d510d6546d5fb07a58cca2b2e07af85c856cc1c35a95388d56c79beb0ff780;
  assign mdsMatrix_4_8 = 255'h596266671008316025e150315e5b1a2c775f211f5f0400137c29b8598c3f9456;
  assign mdsMatrix_4_9 = 254'h28c8e6cf26a4311ba140667f532d5710c828d8651060353c07d211d752c5445e;
  assign mdsMatrix_4_10 = 255'h495bdc653b04aaa85d2f717969d79ea1fd96306ed9780e3cb06ac039e2551ca6;
  assign mdsMatrix_4_11 = 255'h592ce85e733d0117743e74a8931cfcdb3ffeadb6e8c72dd20aaefa9336808d89;
  assign mdsMatrix_5_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_5_1 = 255'h5fa6c8b46e5aba7b95972470ea764714925d44313f1b53dd406fd632aa03f270;
  assign mdsMatrix_5_2 = 254'h2556d914d19ef3613c86aef70026f1b344c3a73400baff1121b131fc4f096b73;
  assign mdsMatrix_5_3 = 253'h1cf7f0a51375f1e8cf506f6c364ca941eb9a1b2d9cea75c7bc91fec9221f5078;
  assign mdsMatrix_5_4 = 252'had2df7322c6552e7d938df0f8943d6b0790c82bffbe24879f82cfb22ab5edfc;
  assign mdsMatrix_5_5 = 255'h50831bf51e2b1147324ed4e6309448bd38ec8374bfa04016ff64039face4993b;
  assign mdsMatrix_5_6 = 254'h221ff1d92e929d542d6cc67918b8d94ccb61cfbd0a6e662003340b3cac8ad19e;
  assign mdsMatrix_5_7 = 255'h4ac6798c23163a468e2ec4822570b9d45b1d12e0396a6428575e70170efd2760;
  assign mdsMatrix_5_8 = 255'h5babbd1d3ac4dbac173857f069694f1532af92f6189ca978070e3adbd5f75f9c;
  assign mdsMatrix_5_9 = 255'h675da5d5bbee23752dabc193ec3629f69864ee522edac81e83d2d21d2ff73c75;
  assign mdsMatrix_5_10 = 253'h10c665c7d1826c227e67d7b297d04e6dcfb3a535e874b4b64cfcf0df0086f17e;
  assign mdsMatrix_5_11 = 255'h5a7b0079258384b69b2dc4dd43c88a47fea5e92ec26e6b216b6f69b35e9dd108;
  assign mdsMatrix_6_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_6_1 = 255'h60ce577c97b8492a537ea020019fd311e0dd6ab57f2c87e5a86673d03b8a473b;
  assign mdsMatrix_6_2 = 255'h513fdbe346e354ba4077c1b3169c950eceafe52a6cebc77554a14429db2eb6a6;
  assign mdsMatrix_6_3 = 254'h345fec3b247480af7de60f0d2634f2ce3ec5247075216f77769ba861654c89eb;
  assign mdsMatrix_6_4 = 254'h35304725247ba29ff75aaa8ce17b094d1d2033fa64cd5794f7e377aa912bac74;
  assign mdsMatrix_6_5 = 255'h60d591856d4addce0e28aace4f3a6f507bc6a5d4e074425a5d6d85a4c108b06d;
  assign mdsMatrix_6_6 = 251'h4fb86d1cec23f0413fc341a5fc380733f2308a5cc8f4e2996565b1061b86ec3;
  assign mdsMatrix_6_7 = 254'h30c453a9a702f6f6345ec4df68b3816f7252949ae2d422d5680e45f0cfbb09fd;
  assign mdsMatrix_6_8 = 255'h404f3190e05291e0c7983072fd9e592d9d7982af2a486ca99f275faef8ad922f;
  assign mdsMatrix_6_9 = 254'h2518565fd0b00187942f3d60bece35ba67c837d25f60bace0a12ade756f937de;
  assign mdsMatrix_6_10 = 254'h333803e5af43589b4ed33e02ae2d5ae4a18d4f76e9a71e602db8dda184f92738;
  assign mdsMatrix_6_11 = 254'h2820aadbab363a17595e127ad383ab3b37237a524496e237e8cabdd5d29ccb9d;
  assign mdsMatrix_7_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_7_1 = 255'h4be9decec1c886731c4878ffce08f4b3d8f3c41bff8a2547f9c88eeeb51d0848;
  assign mdsMatrix_7_2 = 255'h4f8caca36d8cf5d764b60721cb5e34fc389b266dd9a25b06c0fb224afa300a39;
  assign mdsMatrix_7_3 = 254'h23188ae6156e8b9741b36ebb0fe8f0967d039d7e80e0ee9ec5ecf1b3a3c53e29;
  assign mdsMatrix_7_4 = 255'h42c544e7d8d3c27bd86fae416a2558199d1b689e31b722ab143327026b66a913;
  assign mdsMatrix_7_5 = 255'h430493eb4e124d6dac22deb3bcd84fffc9b65ec7edcb6d1fb0ca1098fb300477;
  assign mdsMatrix_7_6 = 255'h6f4bf3f16015046b315a6778267def2b793119dd3d179d3b31cf85630e1e1a3e;
  assign mdsMatrix_7_7 = 255'h5bffb1120939698b70e85cbb363b05595dd6b72dcaf701ee3434449e28191fe7;
  assign mdsMatrix_7_8 = 254'h2fb8ace57c6cfc025ec753217682d98b9923d29a5f17ee6b62677f539f408bad;
  assign mdsMatrix_7_9 = 251'h4e7998449e4458d80d138d3a192ae2e1953a9bf22d8a7ce9c5235ab5c0878b2;
  assign mdsMatrix_7_10 = 255'h5f2a4595db6b02faac74cd0c1a795135fa0ea6043b23912c8e258db0c25c2b4c;
  assign mdsMatrix_7_11 = 255'h5d0f8143e6012aa70ef47d40907b1f9cb13fa234da097515c28e8c8cc6dda221;
  assign mdsMatrix_8_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_8_1 = 255'h61776af8da9af7de54c57d6824e4f25022c3356ec5d638562ed7b69b56f93b91;
  assign mdsMatrix_8_2 = 255'h43a7356e52be15dd3000e21c4930cd7eab0fa9d0c13526fa15a102a94672cfec;
  assign mdsMatrix_8_3 = 255'h6741f227aea7c54a6760407882ba42bf959871c4db06cf93899de6d684a97b2c;
  assign mdsMatrix_8_4 = 255'h46efa8810fab3d85cb98c1a7798b3831c65079ab2cd67733a10b7e849e2b61dd;
  assign mdsMatrix_8_5 = 250'h3f60c2b214a1ff2eca665825b4f72a60922cec2039b11ba8e557397d193a9dd;
  assign mdsMatrix_8_6 = 253'h12da3e1ff4bb3e789f4053907bcab049a8c82f78fe17a70a6eacde05ad52b0dd;
  assign mdsMatrix_8_7 = 255'h4af7a86c4831b9aa86818db808dbb7f714e67c25d037c69dd4bc5ed37c3ac0ac;
  assign mdsMatrix_8_8 = 254'h2f19f9ffef9573dae0cc77a412647e1421b4beb0054f8e38f7be959256063ae3;
  assign mdsMatrix_8_9 = 254'h2175d9b4f4c5dceb4915fb5341cffa4c8751314b4322db9257df88411a11973b;
  assign mdsMatrix_8_10 = 253'h15adc21a39cd5b825b830d798e544c9ea560a6d54bff534f389dd6ebb17281ae;
  assign mdsMatrix_8_11 = 253'h1cfe0c13c7584af76fa2bb280ea42ebc8fa0019f3e242e9c04c928dd9dd8f4e6;
  assign mdsMatrix_9_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_9_1 = 250'h377af5e4bb407cee0e4f6619cbaeedcada0d3579487fe593f5a3508b47c0ca6;
  assign mdsMatrix_9_2 = 250'h384f885809f7506e87a14183cc111071a856a0580600639aaef4f0612b23ba7;
  assign mdsMatrix_9_3 = 254'h28809f42aef9f02adfccdf9df5710ec4c5b3ca70c7c3d98e9ac872c464efeb1e;
  assign mdsMatrix_9_4 = 255'h4df7a9be82cd112d52f5c7fe24a1f7ea58c4989ef33f2d664a4280f53efceac8;
  assign mdsMatrix_9_5 = 254'h35e91169dd1b111e25f64e9ea401c41540973558b7a6470cf7b43d21c6ecf2ab;
  assign mdsMatrix_9_6 = 255'h4cb215d6ef55095d864c310c59218aa9750304810f79a10243d626b94a38d35a;
  assign mdsMatrix_9_7 = 254'h24d527d2a7458bec357db74f40f58542cffce80a75988c92ae46ebd4df86bec7;
  assign mdsMatrix_9_8 = 251'h5deaa9e5b97f1afb6ad32a90a978d4ebcf5d7d63bfe27967570b5d784bae347;
  assign mdsMatrix_9_9 = 254'h28f8f344c77b81027f48b35d34d83eed23e7637dbaa0490c8be5589b71d90de0;
  assign mdsMatrix_9_10 = 255'h5dd88561e7f13e2f3c48db7dc6e778fc7e2a0450e72773b546bc48781a26dd65;
  assign mdsMatrix_9_11 = 255'h481f575764217f1ee0d8efd1a8ce6d4bb68a2a3446d9153955f35a499cfa16f1;
  assign mdsMatrix_10_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_10_1 = 255'h6e6ab51d1b491bcbea525bfd913907b14d0ca75fbfcad69ce24cdf998720ea9b;
  assign mdsMatrix_10_2 = 254'h32a6f47ff8938cb9735274931e703317ae5e69e57a2f1d4ce309066b6ce7f2d4;
  assign mdsMatrix_10_3 = 255'h6dbb072e3ed03b64c9c3e611d10b6137d15330cd9a8f7fe170e6d27b4a1ebeff;
  assign mdsMatrix_10_4 = 255'h596741b70e2e937c784953c59b59133cd20d2557846ee03353988057f591e9f1;
  assign mdsMatrix_10_5 = 255'h605f4f9153af0fbef957e98e05e50ae7e07c11e1614d8808058cfbde7f0853c2;
  assign mdsMatrix_10_6 = 250'h23591d2d63439e9fb4ded98f0bc958ea8c3acba0102067a758f07adc17ac276;
  assign mdsMatrix_10_7 = 255'h6131822482a16e469207b8acbc320a332de4d4fecaa4ad2d05b9bc15501f4277;
  assign mdsMatrix_10_8 = 253'h14ac14d0a6f8415ca08cf1823750df9cbce7e13441fc7dfde6ab1be4a60dc672;
  assign mdsMatrix_10_9 = 253'h1cd34e84b15b0ca87784ea217174d4e1f174ccb9c28739b276d99f8c1cbea495;
  assign mdsMatrix_10_10 = 254'h24129d5196f20968e2a47bb1ef97638a8e14073b6f2ab8ac19461f73f32ba295;
  assign mdsMatrix_10_11 = 251'h7287657f40c1c6ce5c58cf2a912ae96ceb9d43983894749ee8df472c607571a;
  assign mdsMatrix_11_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_11_1 = 254'h3238e8622a95b50b8002e767df40d0cb2fe42415e30ec8d7f9c137680a10a3f0;
  assign mdsMatrix_11_2 = 255'h538fbda9a477d052afc432c204cbd61b3356a71086d92b9330284472ed87373f;
  assign mdsMatrix_11_3 = 251'h58838699a9b73c117c84a91743d12357f0f3a39d041c5d8ebe31727c1c379b1;
  assign mdsMatrix_11_4 = 254'h3b2fa277080e7f5da5906fa7fea831fc4f309a1e1cb8e19c65d48311a1a624ee;
  assign mdsMatrix_11_5 = 250'h2f9cf824a080fcf3fabbcc052c14dd64977c6fd654acb7dd2e094b8e66fc680;
  assign mdsMatrix_11_6 = 254'h2bf93be464b41a4dc24d811b4a4555fe41595ab9cb5ea8510d3264bc3ab8d2d0;
  assign mdsMatrix_11_7 = 254'h27c2870d6a47be9da14647bab5705181af58eabb925d65167531842607d2dd2b;
  assign mdsMatrix_11_8 = 255'h5bdc008008456288d25f8f653bc6bda0347991cf35ac859f6d8a6317f6548d5d;
  assign mdsMatrix_11_9 = 255'h4dac9f379ba7ec5f004d4024bfbc424ac5f91cff26023d7289a6b55fe4bc0d36;
  assign mdsMatrix_11_10 = 254'h26053ab5ae3e394ff5dba98243a7525946ed1a27cd3fa51e3d0fd53914c44ad2;
  assign mdsMatrix_11_11 = 245'h1fb03707093158f2efba7f32200538b2cfc0dfaa76f41614ec4c7a97e0b64c;
  assign mdsMatrix_12_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_12_1 = 254'h372eec7110dfe4e9fc16784b0f8c486c92c98673b323623130fb59650422120a;
  assign mdsMatrix_12_2 = 255'h67c1a3cac236e97d0241cbffe51aea326eda78c2322723afc3e6f9cada292dbc;
  assign mdsMatrix_12_3 = 255'h5b58d527815cb0ee11cce8e3bb5c50d5c302d45365fec1f1e595267732f7718a;
  assign mdsMatrix_12_4 = 255'h5f0aa17442fccb943757e0474c927b88ed735d1adea7673cbb10c3455aa3cb1d;
  assign mdsMatrix_12_5 = 255'h6d84c9e0bbfda7b7bbfb53f787063b5b6054ca3ad5df1a4722cd2e556960094b;
  assign mdsMatrix_12_6 = 254'h20ad06bd9bf864ebdf8b5501bdf18d72b1c90098aefa335370a26b2bbeab2d85;
  assign mdsMatrix_12_7 = 254'h3807777d2415a2ebdc63a77ae67bb0da286888be718d9becd52f5d0f6328f24d;
  assign mdsMatrix_12_8 = 255'h4aadcf9c133a6ed17f03402df159df14aa9511c28f6d733c04cdda893846aa0d;
  assign mdsMatrix_12_9 = 255'h6f7c00f5fc22ce69a71a89526af5a48c4facee40bc913067517b14f40780545d;
  assign mdsMatrix_12_10 = 255'h4cce3572044c293c7d5a9a5a6ee720ec27425a0500028344e4f3fdff03f7705b;
  assign mdsMatrix_12_11 = 255'h4c7d7e025cabfaa4b22618240713441ae7a6e90d8ac279312aa1310ea3affa9a;
  assign mdsMatrix_13_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_13_1 = 255'h601910ff87e0acd410d1a49c916e496daf6d80cae3e3e4ae5dedc52e07f1f0ac;
  assign mdsMatrix_13_2 = 255'h723ab06e52d243aaff16b3f431037a0f1d519f938eb56ab39da6fb66946b30a4;
  assign mdsMatrix_13_3 = 255'h691073097f91e13cf221cacd9f23715c1f49719b0a134f9a96b54fc8a8d09638;
  assign mdsMatrix_13_4 = 253'h113cf1a61f5816dcf76d4471c3081a79d8246915d0814bc5a259600e4cd587ff;
  assign mdsMatrix_13_5 = 252'hd4beacf4171f42473bfe2e9e117d566e3b96a59e164832140e9c4b758ec0c06;
  assign mdsMatrix_13_6 = 255'h5c7304c1c6224c4e9c76ce8dbb4a6e41e68871115e21fb415736d76baa9d5c02;
  assign mdsMatrix_13_7 = 255'h6546ddad1b8ba38d3f21a96df8f0d7a917ffcc610952ac2580203944a34851d8;
  assign mdsMatrix_13_8 = 255'h70dad03d4b5a78b23c09d35a4c3778aad1451440eb14049ced60b5a269bd78e7;
  assign mdsMatrix_13_9 = 255'h521459cd5dd1a38d21a0f0954062f637ec80d87e940242a2b27d9f5c3e6f28c0;
  assign mdsMatrix_13_10 = 255'h5860c31b3265db1f300e7ff70bdacc20090059ed2db7594a9cd93b5e5d20b62d;
  assign mdsMatrix_13_11 = 255'h66da699124d2a311b3f183f2695e619242b26322175a880eda41aeeca5871197;
  assign mdsMatrix_14_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_14_1 = 253'h16eeac223b2e74e5af656b8720ea535bd039ba94aafcceeabac62aa941203d0b;
  assign mdsMatrix_14_2 = 255'h5804aa84719df2f1e67605727eebf7a252bf2ed15c92a2fc54ab6c1cc6ebeb63;
  assign mdsMatrix_14_3 = 255'h51659a8068906d2c5c28b7e06c96ef765802381ca75bbe6c28024188e0a448af;
  assign mdsMatrix_14_4 = 254'h3b87295f0006d6597629a9f39d83121f1e01d8829792cc5504d3060b39b1e1d3;
  assign mdsMatrix_14_5 = 253'h129d9526a82f9f125e3496a712a3bd4667e9e7c0223b81488b01159f85c3d4f3;
  assign mdsMatrix_14_6 = 254'h3c7a5b68f2095b7735f86ceb143ff86c342ea1338ad2c633484f14afc2a42219;
  assign mdsMatrix_14_7 = 250'h3a0c6428ac63e7a5a5f88c4c9587efdcaad9b295b0258134efcd851321a8870;
  assign mdsMatrix_14_8 = 253'h1d06e5fe365487997fd7bc412cbd8d53420c2f5c7decda096fc8236882c36ba5;
  assign mdsMatrix_14_9 = 252'hc54789084e9ea5359a608282b64b6a59bde4fcbb88f0cd244257df313710565;
  assign mdsMatrix_14_10 = 251'h74e43b8c22d1635c7beb16caa133d5d7dc69ac16431a67d47528a8c2fd8649b;
  assign mdsMatrix_14_11 = 253'h1c3d8668c3dcc02d0647059b4ff08e076967845a6779e4f93b44aee5b7df12e2;
  assign mdsMatrix_15_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_15_1 = 254'h3cc66d55fdd590482137c25652c090496af332539989884de5dd41a6e7dc635c;
  assign mdsMatrix_15_2 = 255'h711b196a75cf35230ea37237173e2e55816eac1308c90f0bab5fddb3995eb847;
  assign mdsMatrix_15_3 = 253'h1f87106d80fd41937fe5f7f9158858f80f2fcec7abda7ebdb72f8d3d36706e66;
  assign mdsMatrix_15_4 = 253'h1cf308b5463ec249f6f1ec6dc8303d0271e17c6ae133496f3915f9f87df7dfd0;
  assign mdsMatrix_15_5 = 252'hca0d70c556b411055a8f8f3042e95545b3698b0d49bee0857b870a0ef99e0e4;
  assign mdsMatrix_15_6 = 254'h2302a76e60ff1bf346c90fd1aaa9233d6b843ad6e50b724c5689e56c392fb195;
  assign mdsMatrix_15_7 = 254'h25ef1688dda223ada5932f0f63d896aa2216508b955fd279f893cc9ba8948c57;
  assign mdsMatrix_15_8 = 251'h6532dfeda6ec9fd6a2b283cd6b2f6bf636f3ceb11dfeb1d27998a141029a6aa;
  assign mdsMatrix_15_9 = 255'h4cc2db604cf033d747b45ed206aadea6c7b8ddcc42bdb38f14999f62d92b9e9b;
  assign mdsMatrix_15_10 = 255'h72ea8f97cf887e0c023e2060923c7b984f212e4e80aa16053c18d46469bf24d3;
  assign mdsMatrix_15_11 = 253'h1373d2377b57277ca7aa4d16c3a676712f94b56483614292ea3c64c6d24b5c77;
  assign mdsMatrix_16_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_16_1 = 255'h64e2146eaa916c6b51c3c36a61a98cd360b24ca61c9f89c29c62f6f855ad5c54;
  assign mdsMatrix_16_2 = 253'h1f07aaab7180f2d9b189f6b5b27e6f2530e38f09df90589404b493d60be17553;
  assign mdsMatrix_16_3 = 255'h44868e9d140e507f8d4c972b928e9eeabc88951a5f1091228dba9ba1b3c2b6a1;
  assign mdsMatrix_16_4 = 254'h3a55a1722ac52e623fac5aee85df711e911c781e4fc7225d48d5d1ad49f3e825;
  assign mdsMatrix_16_5 = 254'h3cbc6dcb970c1776e2ae5e84bc27503494a7292d00213e66d5f8753a40c45f31;
  assign mdsMatrix_16_6 = 252'h9208d41936a8b6a769e9ad83fb8aa09286395b3a4b37b0413b50327f1725b89;
  assign mdsMatrix_16_7 = 254'h2688605373af50b6e40c625aaca0bf6bbd53370406116faa247a31de08b6dd5e;
  assign mdsMatrix_16_8 = 253'h14547ea6932c763817dada904b8ff1b0a4c641ec20f3539b8511d35cf1d8ec44;
  assign mdsMatrix_16_9 = 254'h2feb901a2e7218a605ba88404cd1a13ef4b83c50f40c4baf007543133d0768f7;
  assign mdsMatrix_16_10 = 254'h28bf58f510becbd771440bc3f6b430053bab2793bef12afd69667570f2dcbc61;
  assign mdsMatrix_16_11 = 254'h227a62d3b81950b968890db1fde084e2badff0e7c15dbf53a53e3734797a33cb;
  assign mdsMatrix_17_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_17_1 = 255'h4b92b931108e2892a3fbcea26839bd544ea4a83954a0f80279c0ad1b510c319d;
  assign mdsMatrix_17_2 = 255'h41f95d89dfe0ec1185fd386dc840d28d613a869a12a47056b3ba9620319ad627;
  assign mdsMatrix_17_3 = 254'h26cccb0cd28c8b8292aea871fdca9eb807949329b607eb9afb86c50d1b262bed;
  assign mdsMatrix_17_4 = 254'h374803f6710c998df325f772773220972016636412d3d05d8a9d778b14a15e00;
  assign mdsMatrix_17_5 = 255'h4703debf82b07f58b8d4a9f5c6547fdf3f3039e7163f813ebac320df53170c85;
  assign mdsMatrix_17_6 = 252'he86ad3b151041d9999b98894c5efbbeb000419b35907fb5928183e5b65350d4;
  assign mdsMatrix_17_7 = 254'h252d65bcbb52cb883d980b80d5f321b3009a64e860bb0b2c6a62a7860626e2d7;
  assign mdsMatrix_17_8 = 255'h4c0b8b34eb5374c2f151c0912a099f7b6b0f35be0634141256a0965769ede152;
  assign mdsMatrix_17_9 = 255'h6985542992b8b652bfff64b282fac988929ca5b4561865b7723f4efc2263de2e;
  assign mdsMatrix_17_10 = 253'h1f9569e3f5201e9960c9f0647b4f55d24d807e8337539e84914da50fe6b49971;
  assign mdsMatrix_17_11 = 255'h6abbd7511ffebae2239735952021d5e31539526f8d03ad932cdd9e0f7f333575;
  assign mdsMatrix_18_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_18_1 = 255'h62c61b9229f3b0e37510ef1c72ac36ede2309cc7fe2be3d4f84481cef8d8d83e;
  assign mdsMatrix_18_2 = 254'h2312fa1e8bf66ea8aea0da7581cc1e5061aa23ea1f25a3379e0e4206235539bf;
  assign mdsMatrix_18_3 = 255'h5c7ca826a71aa52838ae7164e41f244aa5a7f179f68ba20c078106c4e1fcd5f6;
  assign mdsMatrix_18_4 = 253'h146e06c7ffa98c2bddc9fac5fe08d6012e8121a800b609d21685321e7f40b85f;
  assign mdsMatrix_18_5 = 252'hd792ba8744347477927e19d9b0a01514915a4698fc7db69e5f8f06a735bb96c;
  assign mdsMatrix_18_6 = 252'hda39d4d1a6dc7b4a6845f0fa9a778b37f14a8c42fe345e17ac074cf8cc705b9;
  assign mdsMatrix_18_7 = 255'h46a86873e7de2109aeaa764623e3cbcb40186c0c72960f496f9fb9452296815f;
  assign mdsMatrix_18_8 = 255'h527193335f7779c86b99245ad5d69e47ac8d957f7c286843ed84456b54fb5f9f;
  assign mdsMatrix_18_9 = 253'h1c0a6cfc9cbeeef53a09a76620e55a8bb6f4843a644e10083e82a64a44b2382d;
  assign mdsMatrix_18_10 = 253'h121a45e7bb27cf86e3e6eac5febe26a001c4ae26fd3534f3d41db10c64a2f76c;
  assign mdsMatrix_18_11 = 254'h2b7dba70dd1afccf1b9c6be2fe30413a3106a2dab5f9e465b345ed9d5b26505e;
  assign mdsMatrix_19_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_19_1 = 254'h36f2b9cf006cdf1b45a0cfd8307e5a7e0d6e6c82aaf4e9156b62466bc35386ac;
  assign mdsMatrix_19_2 = 252'hbef6b1f5ba46332f5df9528bded15a06e8535fc2ed2dd134848279a98051b9a;
  assign mdsMatrix_19_3 = 254'h3ea6a553d0011039081601be8b6086ffd9001cc8660e1f04a62aaef29e6a0b9c;
  assign mdsMatrix_19_4 = 254'h29846c1c3171ade0b52700db82f5664650864776f5f65af0295885435f9a19fe;
  assign mdsMatrix_19_5 = 253'h18f2aefebd03954b21b177a3ee4d07a3e525b72772029e66becb09f0f9e7a4e6;
  assign mdsMatrix_19_6 = 255'h411a0005a1c697860a66e49727e4fb1797101076c6d025ecd77ca3d0ea374af1;
  assign mdsMatrix_19_7 = 255'h532294cb1ee44d1e092eb02f58bbffe771e9b373f7b6781dda7f42357f238ae6;
  assign mdsMatrix_19_8 = 255'h5d3f09996c229b26e891e683f79f8131615d6168141ef93c8de08c240cb847b0;
  assign mdsMatrix_19_9 = 254'h29a790dab3d55e5eb7e07585daca3e3b6a146c904e8efe8f3f8268bb2c5bc5cb;
  assign mdsMatrix_19_10 = 255'h599078fbcd661b1f5c60d9150e46033b85a860b8bd28c7933fa52de2d743ced2;
  assign mdsMatrix_19_11 = 252'h94673f10b2f65489ac1a815cdf33cea76ab964a323ede6180cdb4998c86d0df;
  assign mdsMatrix_20_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_20_1 = 255'h67d16e26dbcf8e8dc59a1a14eac79024e2297f58ef3895f2a53fa038466187b2;
  assign mdsMatrix_20_2 = 254'h3407007e6179e15b976e114cbc44fa0969508bf1bff05b917a25e59778cfcfb6;
  assign mdsMatrix_20_3 = 254'h2ac4344149e8a0c2b74c52e33e2546ecfdc3f143450ccede6a3ba7d79419504d;
  assign mdsMatrix_20_4 = 255'h4ae4007e4dae2951ac771d42b3fe7a8c76739bb3396dc1b6b491f2e777171fe6;
  assign mdsMatrix_20_5 = 255'h45ed2ebffbcfcfed7100f0f79f169690383d79d7ca0c2e43e37b38455b065125;
  assign mdsMatrix_20_6 = 255'h6160a3a75203f7b110260c667e374241a9cfab6f94ae5fb03987f6162cf418ef;
  assign mdsMatrix_20_7 = 255'h62c7c1d136e3b1cad2acf4e5fe11fddd449a56c6483d44ae0dd0c23150c445c4;
  assign mdsMatrix_20_8 = 253'h164b09c1088bb7c7c3f8e8cf1f31f08ffd6ed49e6afc6237f3cc955d5119f71c;
  assign mdsMatrix_20_9 = 251'h5651a8583e9cc008e06a2ee78de60bca503d37f5a8475b2028f888866566a97;
  assign mdsMatrix_20_10 = 253'h1d142e92b853d3453ef70bc433a144a24e1fe6297a27ecc864b0c9661f38b24d;
  assign mdsMatrix_20_11 = 254'h291630e1c304b295751db4a7264c513ab45bf2acbf19c781c6eae16f02a95f9b;
  assign mdsMatrix_21_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_21_1 = 255'h4643ada1732013335de9ea52412b52539b992c6649de0779969626ccaeb20881;
  assign mdsMatrix_21_2 = 255'h4cadb5edecd50b6e43c7b3d33d8d49fb3a37ee1f480fb5987a3690e69f2e8a9c;
  assign mdsMatrix_21_3 = 255'h53cd0947ef252cdc69c8236b5d9cf62f8d95f982381df022a22723fe2863e5d5;
  assign mdsMatrix_21_4 = 253'h1d89372084d3e8df48bf3f5340b288eec67df9988bb461ee00fd665f6088a7ce;
  assign mdsMatrix_21_5 = 253'h14ccc00196732c0ba859d999ba170165775d5361af6b4c3e720fb55fae0c2f7b;
  assign mdsMatrix_21_6 = 253'h1fbcf3b07c02ab41426043b25647314321bca92751b441005a4e37c7fbbcb44b;
  assign mdsMatrix_21_7 = 254'h25e2634105db92126b6a54da63892776206d3f30183fc148550c5d5cda2b6d24;
  assign mdsMatrix_21_8 = 251'h498aff10d87e8ab03bf4f914c5737b254a9c6b7ffdebdf23330fdaad3718666;
  assign mdsMatrix_21_9 = 254'h27f36ea3d97d69858789d999fdc4a82723a7e1aae297c2dab56b7497b425c0f6;
  assign mdsMatrix_21_10 = 252'h914b4e0cb46e9ea5ac7acccd390dd9b1dcab9df0704a70cab3b6a63e1901a05;
  assign mdsMatrix_21_11 = 255'h653276b852f574742654a66d66622f98660dcbe26ede67cfe964d13d145b61a5;
  assign mdsMatrix_22_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_22_1 = 254'h28e361ca88cfa602c6263366aa0e381659bb8ae70f556ad866056ef60e199dfb;
  assign mdsMatrix_22_2 = 255'h6cc6906f4aeb828df62f7481e0baf9d677eed9f36312636f8d3c96889d3d4a78;
  assign mdsMatrix_22_3 = 255'h6dfd9c53363835cc88bd0c938d40b3c968e2a9be80bffd7034d9809eb095e062;
  assign mdsMatrix_22_4 = 251'h790662d205f5fdc1733978aeccdb1e314eb12eb089d9eddaf735e2f451f368b;
  assign mdsMatrix_22_5 = 251'h71ceacc24e9f9b37fa2b4ca5cde7aebd4995d8602393706abb2501812c6ac4f;
  assign mdsMatrix_22_6 = 255'h4d3c180afb7192a4da13ac4db67c0e1adaee25064aa50d123999ac3977c619b7;
  assign mdsMatrix_22_7 = 255'h7249259500cc4a9542e05b7a69b7759a700f2a0464c427dbc4bf60428d5a3916;
  assign mdsMatrix_22_8 = 253'h1b5f4cfec1b35474e0db44e60299d47a9ee82c65ac4618b4c919eda216bdcee7;
  assign mdsMatrix_22_9 = 253'h18fe0153c0c594dfed29815129f5274b98108d3ff9b3efb842517aa452a7663c;
  assign mdsMatrix_22_10 = 255'h6dce8b7747aec312058de88431a957cb028b254b1a7f85de2d364c40d0ac0cd8;
  assign mdsMatrix_22_11 = 255'h62ec82913584dc414bb87e4439c2975b26f4a06f11c117c54fc925be3f548693;
  assign mdsMatrix_23_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_23_1 = 255'h550f610ac51caa9d15301247002dfc92a878e614505fa680c389ba5c0931894b;
  assign mdsMatrix_23_2 = 253'h19c7a97d7a9c30f78c051e6c9419212ced9f5fe00e71d421f34aa97396c18deb;
  assign mdsMatrix_23_3 = 254'h304354f6db1fcfac69f95a05055f291ae2ea554795336cca33b2f0f3e8db1197;
  assign mdsMatrix_23_4 = 255'h56dc4ca87f58860d70d167b0e273f0ff358903debcde9be0219588a2eb67bfcf;
  assign mdsMatrix_23_5 = 255'h6fcabb67462a670fbb75e9fdb583f72cf99159be4497fa517f8b1e095171efeb;
  assign mdsMatrix_23_6 = 255'h5a7a60c7e07bdbbb426e0d86b94489d30cab471528bfdbf565b07789a4c03075;
  assign mdsMatrix_23_7 = 255'h4167dc9e12bea1506c65864b66620c7159435d0e4e9e2d8207b4bb7dea6e9826;
  assign mdsMatrix_23_8 = 250'h3841263b2efe68f3e82ff7c243ae948c82867d6a642bd8d6d4e1f34d18f76a8;
  assign mdsMatrix_23_9 = 254'h29ff6c3b22c584995cea3f7a71a67922deb538b6a844e4c9b33634861de83cff;
  assign mdsMatrix_23_10 = 252'he91b44a72c2531737aead8fc004362503047c030b011c65d3eee0461468ada8;
  assign mdsMatrix_23_11 = 255'h500be8fe5300dfb084b504f7ddda6c96b71a33e10c1be04aa6bee52e79f9972f;
  assign mdsMatrix_24_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_24_1 = 254'h3068f6369ec8d2bf0e19d8ce8a706aa9502f79b455f28a0f91f8d058240585d1;
  assign mdsMatrix_24_2 = 255'h59702a9bdaea4365f2b619467bdc512c8d2f450a5f4ad9ac34c71403369e7d99;
  assign mdsMatrix_24_3 = 255'h5dfaa3314124269bcb6a3ec5e1100a635807ab527886a202ed633e75c5310b85;
  assign mdsMatrix_24_4 = 255'h5b1defddf3c3068c47ec7ac884b61d0a433c43a4ed3d7e65b267fe8e6f8c0ce9;
  assign mdsMatrix_24_5 = 254'h33fffff19c0e9422a908dda78783f780749d529fd79e9dc0d44a2cbe2c334e5b;
  assign mdsMatrix_24_6 = 255'h6d01cd556b963341af3e45f3e0fb3d3a2ec1c4f5add7ea8240518d07ddfa9657;
  assign mdsMatrix_24_7 = 255'h6c6c5cc11245ca4903ed1f811b6e4adda886f3dc700a6ac18ca45fd0deb43504;
  assign mdsMatrix_24_8 = 255'h5fc72d21bac0c95f505e79d7dc97063778bff2580d25435681e2c1fc53a6d46d;
  assign mdsMatrix_24_9 = 255'h66a28682b30a6760464a76b438b22c4a8629ccca270a2a94a82634ab1870914f;
  assign mdsMatrix_24_10 = 255'h6dfe1f14c3770f2babf18729e7db07dc9c7154c0848d337d849997d18541abf4;
  assign mdsMatrix_24_11 = 254'h387cf23f1195dac28a30473e5f4372410d3d2ccec747b93b37f2f55595f7fc60;
  assign mdsMatrix_25_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_25_1 = 254'h250deda6a2e431c4f6601cb52f96cc858c5f015ed309408cd6023af2e4067ead;
  assign mdsMatrix_25_2 = 255'h629c4fe76b2cdc07fe03d9a55b6e0471c49e01de13a591013db8a15d704b27c1;
  assign mdsMatrix_25_3 = 255'h423d01a5ad424cb7792e09b4d187db705bc69b62000a81a8be0872064d033e8b;
  assign mdsMatrix_25_4 = 255'h709b09e5fa990bdf6fe18b25dfe6d7276f4812e5fa79bcd6696f580b850e3700;
  assign mdsMatrix_25_5 = 254'h318123df6d69237e16e27e51aebea8a38c0c89e38ae9881fbe63df72348b54c7;
  assign mdsMatrix_25_6 = 254'h3708328818cd4e176e0cd927d658a2ce39eed921437c20f2a635d60acebedcca;
  assign mdsMatrix_25_7 = 251'h4264f88e7049d77537b1d2b847efda3c6e58d1638db8ba3d6a1c05897b8dd22;
  assign mdsMatrix_25_8 = 255'h4ebc194b978b975b0ad75fc67342f6dc7f613771e5bab1ed321edd6efb9b1c6d;
  assign mdsMatrix_25_9 = 255'h51fc091a9be822727f2177c530328b8ac8fdb2126e52de20fbf1a55464f2f35f;
  assign mdsMatrix_25_10 = 255'h491390485b1fc91b6a7e00da41a0e1cb98ade02bbc2bba0cb44e96167211da44;
  assign mdsMatrix_25_11 = 254'h2bacecc7228e36ecf4452a771b2948f161896c73c272e425eeb8032b3825b7c5;
  assign mdsMatrix_26_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_26_1 = 255'h4e0b5a8f8850a9994cdee0da4be6980d401a7a9015ea7ff1456c3ad90b3084fa;
  assign mdsMatrix_26_2 = 255'h6fedd284f52b1dc752a09915946bd84f180d91d2005de3bb0c1071a4ebd2a3cb;
  assign mdsMatrix_26_3 = 254'h25ad9cd40270aa89b03fb620db36f5a3a1fde9026a3d13f52e1117d44db7e7d0;
  assign mdsMatrix_26_4 = 254'h26a967780ce80470d9201cbfeeb755dd8e4430d95d11338da24c895308962ac7;
  assign mdsMatrix_26_5 = 250'h2cf78e96ec5f64e957c683ebbef314b0f04aba42bba5556f9cd901b91497aa5;
  assign mdsMatrix_26_6 = 246'h3bc2ab704d82d5317970313ff264dadb9536ba19922837884906642342fd3e;
  assign mdsMatrix_26_7 = 255'h59fc6f552ecef8bca10bd7986090e48aba1d17c595a5d716db39eac9352ba56e;
  assign mdsMatrix_26_8 = 255'h54513124a33483cf03e0e7c932d4699c5e2d8f4d39d165448230d517e9c271a7;
  assign mdsMatrix_26_9 = 255'h6d48b72b1a6aef6dca175128fcf48f26334fafec5a1172871959fbfae4eba4a5;
  assign mdsMatrix_26_10 = 255'h6f09b8f0e55495dcff7e182a1977cd0f90055bcff1ccf1e6adbf75f80c497763;
  assign mdsMatrix_26_11 = 254'h28ce140519d716bc20a7e7c1c6ce647ddc78ce84539d7dbfd97b6cc4ec52b110;
  assign mdsMatrix_27_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_27_1 = 255'h6050a23b7157afbf43a8a4b04b2709f0ca58e725d1a2eb9949af01f2407cac1a;
  assign mdsMatrix_27_2 = 254'h2bc009def64b9e2fbec12f554e2a56b90848e60094829364a9c9d4cea69b296b;
  assign mdsMatrix_27_3 = 255'h40c3ff0e65a6711e6bea0c1ddb4e772e589f2e1f1af7ad73f4fff7a2f25121c0;
  assign mdsMatrix_27_4 = 254'h366ca21156ce6635550731b9b5078541f9b3eab9204ed8dc481501fae5e7a17c;
  assign mdsMatrix_27_5 = 255'h52a7bb3d447a2f45bfceca549bf657b4009652093d19eef9c0bf568ed222d3cc;
  assign mdsMatrix_27_6 = 254'h3153ca176638759e4c8b3d794e07aac63874b49df05e4bdc07aebe5e81183a43;
  assign mdsMatrix_27_7 = 252'hddc79831082eb0a670340e419f6f8cc957f523393b25db4b5354368a5e2a9ba;
  assign mdsMatrix_27_8 = 253'h192e7cff71bb90785b45720decf8fe29ae1deffde113489ea0cb5e923f962c9b;
  assign mdsMatrix_27_9 = 254'h320476b1321ead1044ea706654dcaa503a757e63f181180ee89cc9e2012aefab;
  assign mdsMatrix_27_10 = 254'h2f11c40eb8b01e558b8ce9ee467dd869ebf50d262c324710786ea248a02d6bb8;
  assign mdsMatrix_27_11 = 255'h578b97d3717f38b152414890a7a2017cb353e187091d85c9661d933fe5617d5d;
  assign mdsMatrix_28_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_28_1 = 252'h9c14cbb38c17ea0b915a53554b9908bf774fa340aadb091e1d15540fc18bb47;
  assign mdsMatrix_28_2 = 254'h221c4a13163f2ca5b7c76e66560f29078358615881aaa84d8d1ba261f1d21a7c;
  assign mdsMatrix_28_3 = 255'h6ce5e1a02ff6b25fcc2c4fc07d3a2e27ea215a12d21279a376eef41f4d27d667;
  assign mdsMatrix_28_4 = 253'h1a94c185c124a28e6e7b9f4587ecc09dc9ccd1d6d82aee26dafe99429147f51a;
  assign mdsMatrix_28_5 = 254'h2fff43c8a48c3635eff806bada4a5cd2ca5de2cf6b8064c26cc9edef5046e18c;
  assign mdsMatrix_28_6 = 255'h54b46107fccc85285e6329808361ed1365f6ab9b93120dd6bceccef08db97707;
  assign mdsMatrix_28_7 = 254'h3bb4e7c382bd17926511eafd24e49488c9be39b3e8d555b71963c9fa025fbe31;
  assign mdsMatrix_28_8 = 253'h15cae9bcc60fd9c715c8dc80c15b8058e52bb4ccf1f599dc8083afb13bb66a97;
  assign mdsMatrix_28_9 = 255'h6fa1a1f593aa72fea847178826737a1b726a5212f59ffb7a32d781a2de0975ec;
  assign mdsMatrix_28_10 = 255'h590a88d317be6e47b0aa0967e8ae8fd95cad3215b9f21349def895dfa5500151;
  assign mdsMatrix_28_11 = 248'hc82c37d3215175d9a7073b3beb5bef3ff46433c1a4170d4019d5192b2f8e7f;
  assign mdsMatrix_29_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_29_1 = 252'h8368399dc6b812443dfe0ecae2365a76e04730307ce41b0e55451200100aa75;
  assign mdsMatrix_29_2 = 254'h3e25653239fa221f4ff80f1965d868cf98df03acdf997e92bbbd21e24510fc63;
  assign mdsMatrix_29_3 = 255'h6da6ba7594bb469275126f4c2ace2c9a608308471fe38b82c528d8844134b786;
  assign mdsMatrix_29_4 = 255'h6b7ab203203371d718b35c3768b513202ebb5a84bb4d5915895306517e5c4a28;
  assign mdsMatrix_29_5 = 255'h516a1330845fd881ed3a3077769ffcbcbb49b5f03f3bdbeb90b87246128a6cc4;
  assign mdsMatrix_29_6 = 254'h21a1ad2b76b393ef9b64681c9c43b394aeec7a08189d6c73a46d9a108f150233;
  assign mdsMatrix_29_7 = 255'h6e0b186f0ee722c64511660572dce8239193bde8e60ed269ea1fa31d090503df;
  assign mdsMatrix_29_8 = 253'h123b1d2f5d3337dc2175c1ce31a6ea5616f3db7eb61ee95f85a86a3884cbe079;
  assign mdsMatrix_29_9 = 255'h4c95352b7e8459a7e7951504a33c34fc171f6a9dd8b96c4da6e135c487488d15;
  assign mdsMatrix_29_10 = 254'h230e5bbbc78970513d557677b33b77630307138aac731bf420ad7c2e858884f8;
  assign mdsMatrix_29_11 = 253'h13e632cfbfb03528a859222540ac883ccd4b2305c94913c1ac8ba64d3536dd23;
  assign mdsMatrix_30_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_30_1 = 255'h41e5b0e7671b34aaebbe34c38e4a524ea1cc1785834ed9e324ffb79224a96ba9;
  assign mdsMatrix_30_2 = 254'h3d6250d5ff75268d3a01f17de4c275caacfcf46e033274a68d4c51a302a15f0d;
  assign mdsMatrix_30_3 = 255'h5da3c9bac0c201dc79544e6ff6a6606dd86c9dd21e38e8e011e9fd6cbc56a509;
  assign mdsMatrix_30_4 = 254'h3cefcf7d2d735fe6042806fb935d8b06d9e86d670fbaff3ad42af5bc97b22ce3;
  assign mdsMatrix_30_5 = 253'h1b378a11385f1ef97424a21f00aa478608d33eb00beb74245394442ffb946311;
  assign mdsMatrix_30_6 = 252'hb6c30a48f1dab990e5dcec0eb0b96fd6dbf4788f0be66db94679cbb9396af2e;
  assign mdsMatrix_30_7 = 249'h1266134f47176fff8d5e91b15c5d6b921ea987368de4afe3151062e199559f5;
  assign mdsMatrix_30_8 = 255'h469f186293f162d0e7fc3c7041bdfeedfeb907ef9b16fc7d9720be6d38e5ff41;
  assign mdsMatrix_30_9 = 253'h1a32fb863941dbcc57bf2482d53b915c234fa4f6b5866a51762d5024b5a84501;
  assign mdsMatrix_30_10 = 255'h4f57675408f3722079a862078170cc6790334666992424bc32f75aa0e062ffeb;
  assign mdsMatrix_30_11 = 253'h1fa7132bcfce030f70d61f1b4b5a53abd2670767b13875d1238da0362b4ec1d2;
  assign mdsMatrix_31_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_31_1 = 253'h12bfcd612bf63880432e7f48ddbdd6b45a069e4b5182fbfaea718a4688006c72;
  assign mdsMatrix_31_2 = 255'h4dad2af68fcfe11ae03555b1aa5d179f4c17c414b7f0d48689e05efeca121394;
  assign mdsMatrix_31_3 = 255'h609b61f0df7eb8e4b07495627433a51f90b54b89574f06abdee8be377fa2d944;
  assign mdsMatrix_31_4 = 255'h4bce47cc734589ef6424a4f6f2e12baf761c7f462d968105ac9bec5c2c78af8c;
  assign mdsMatrix_31_5 = 251'h48cf7c16fbed0d3faa29bbd8ad103b0461bca08d3250f53c75007cfc61f0655;
  assign mdsMatrix_31_6 = 253'h1646776fea7f7f097398eaa07785a5658e23d5ea15af9aa46a7c9f9d26a9b2b2;
  assign mdsMatrix_31_7 = 254'h216d1e4e86ecc851fb9ff9822c65a9b02ab8f2a7cee5c708197a3d345d0f39d0;
  assign mdsMatrix_31_8 = 254'h3f1a149520f6bb188c54f016592812e9a2760413806d04b3d57dcbfab30c8290;
  assign mdsMatrix_31_9 = 254'h28e4106ccd4bc81ae77fa90502157f54a98e9db447fa9891f4b90f47106a9745;
  assign mdsMatrix_31_10 = 255'h6ebf90917892f98dc848ef8c853f06a53560db2a0d62d2b9f45b3b7055c30e18;
  assign mdsMatrix_31_11 = 255'h58a2aac3ec8bdbb10936701f50bacaed25a2765524d0fb57f5a04e170a929778;
  assign mdsMatrix_32_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_32_1 = 255'h713244a23e393f57e389e5ab110c76d47fe36adb2b4bbb0f21d682a11956aec1;
  assign mdsMatrix_32_2 = 254'h27ddc08c1ea3e620771e4f923181e19b59c5150c909914d6798cb533fc003dfa;
  assign mdsMatrix_32_3 = 255'h73ec4d4fff2b5775fce1a7b26b51961743e53788860187517c47777b75e49b8f;
  assign mdsMatrix_32_4 = 254'h20fbc29d7c81da9edb745c4c077a940b28c7f3c4350f16d2345533bbe204c1c7;
  assign mdsMatrix_32_5 = 254'h3bd1c105fd75305ac69c8c9a4285ca94e0049596d1159f8ad18dbdcb5a459ee4;
  assign mdsMatrix_32_6 = 252'h93f25f45f1539c933151d4278f40cbe8413ed840d6b0033d28eb1c2e5424910;
  assign mdsMatrix_32_7 = 254'h3555df9411982cc50dd421d172a3e6f9cfbfcba4d6fb2fb23a88f146f9466652;
  assign mdsMatrix_32_8 = 254'h2079a2f649ec32017682cc29225c08337b850c3e5cfb46b12dfc041e481bdd91;
  assign mdsMatrix_32_9 = 253'h184eb7a2e6862549978fd52eedefb8ab680eafe72fbb1444951c812955d9d2c4;
  assign mdsMatrix_32_10 = 254'h32e69d77e2d032fc5d5a6b4ef7c1d9c2c9121532a4036bd3dfd6fadf949c8bbc;
  assign mdsMatrix_32_11 = 254'h293ea9ef270939b6b4af74168268b62e7c8c90ac220f8d366465c749117b7669;
  assign mdsMatrix_33_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_33_1 = 253'h13a8617340d1bed2d3943fdda7095ba035bb01a260e150862e1ed92131dbc862;
  assign mdsMatrix_33_2 = 255'h44902f048498155f94ecc84216a5832221adce0c8a5bdc90e1745bbcb89c878f;
  assign mdsMatrix_33_3 = 255'h506340152e63c8492c4b26f06b67f90ffe577a13584d3a0a989551ba2f8d98c3;
  assign mdsMatrix_33_4 = 254'h2f5db7ac382588a8ae7f7d5c963be6e58ae68957d92f1404348951e1a6bd047d;
  assign mdsMatrix_33_5 = 255'h4186b03e4dd03340ae67ce0e59c6cb33888419893f9c03994cd614f8abfd93a5;
  assign mdsMatrix_33_6 = 252'hc6eb70dcfbf89ffa665596cdc3df431c3ed1a935746255893c65f02c9deb7de;
  assign mdsMatrix_33_7 = 253'h129bc6708bd74abf7b01240c12510600e6333a983d32d827b2101285e19ea1bd;
  assign mdsMatrix_33_8 = 255'h6f1b3c08ce8feea1dc8141db06073578835739f4b7574a300acb4fc96098f750;
  assign mdsMatrix_33_9 = 254'h2415ac39d1a14a6c03a4f7468b4376214a7d80b156744fe67ca4206b2613715e;
  assign mdsMatrix_33_10 = 254'h35b16cc8f104cf78cea3c3fd80a5db81c4a7817616d436240efeac3c58af042f;
  assign mdsMatrix_33_11 = 255'h4a5d2e20ecd88eb1fb23f002c506d8900b1eec7484122a8ce6499c09e4a6b323;
  assign mdsMatrix_34_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_34_1 = 254'h21a486261ac2431f23858de3cd00f0df30bc42dff00da9099c9c803f2c16456c;
  assign mdsMatrix_34_2 = 255'h4da7c5a96b15c41224789c3a9938316147c5ca07097338429172dc67e2044223;
  assign mdsMatrix_34_3 = 251'h645ef104d9b2bcbee8bdfc16a399c9d5f01fb31d6cb5515fb414d03dd2121e1;
  assign mdsMatrix_34_4 = 255'h5637c34c57d7be7ef4a65139776c350fa3a6fadcedb34c898187096eacfd3dd6;
  assign mdsMatrix_34_5 = 255'h63ba4a4c6af3f4e5cb6c9b5fdc4eb7f86b0d0f09f00fed8a2934140d744c8bf9;
  assign mdsMatrix_34_6 = 253'h1b506eb61ffee5e016852db08a575fc77118f0eb15e84661529f5a0fba4723e1;
  assign mdsMatrix_34_7 = 255'h6f082bf247ced25ab8226dfb3aa540794057e112ad37812e99e5ad4d79eaae47;
  assign mdsMatrix_34_8 = 250'h388be1d6d58130225b4c8212d39621530f57166a61563cf003ad2476ef2b9a3;
  assign mdsMatrix_34_9 = 255'h501035c1ea53079c362b9e2e788f2b0f7108aa7d65013772751e291ce8b86557;
  assign mdsMatrix_34_10 = 254'h237d27720223e292b4acd87b23e8015328bb9d7ce6c537eccc850c6b2757a760;
  assign mdsMatrix_34_11 = 255'h47c94a7c976bd517edbf9e5cb8052137cb4b68498c44dfa2d32b5e7ab42eabc2;
  assign mdsMatrix_35_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_35_1 = 255'h518ea87fc099c72511cde2b10bfab81687146459cd407dfbf4088b944f92283c;
  assign mdsMatrix_35_2 = 253'h13c7d3d7fc640c4b41c58637ba2b207e354ff3da364f07b8ed6bf2d6c4f5c269;
  assign mdsMatrix_35_3 = 254'h37966407043ff29fb73e9534889df60ae4b6e3f9e93f7134c80ab5eaed848c2e;
  assign mdsMatrix_35_4 = 255'h6ade9262ab99d7f9aa719b8befbf0455a8a48e0adb3f6a6bfe4f86c3cb794787;
  assign mdsMatrix_35_5 = 254'h227b48c9006287dff979ba83356999c684e421803488df4f7da4e358507b98f0;
  assign mdsMatrix_35_6 = 251'h74d8746b67c7523484f9e58df598596d5a81532e5c57860d216700e2b543073;
  assign mdsMatrix_35_7 = 253'h10a777db5f05e93dd91c443b5593354e3b793abcc409a15a9d613273aa773c77;
  assign mdsMatrix_35_8 = 251'h49101874a1d837d51524e5d6b5394cc5d839921eb339d1688820641f748242f;
  assign mdsMatrix_35_9 = 254'h3e2e333dc86f862e4d28c90230d07b256075585f05706b716c5b1a42d1c979fd;
  assign mdsMatrix_35_10 = 252'h90c55dfcd2ce3a9335981d035f6ae68fa829f5221a5c9753594f499d20e6cdb;
  assign mdsMatrix_35_11 = 252'hf393c1463b5207067e4d520224804e298622fb8eb2a677ba6ad13e5bad3358f;
  assign mdsMatrix_36_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_36_1 = 255'h6070359742f18b0fd7b7a294093ff05219703f0460fc21dae7ab2d337e83ed1d;
  assign mdsMatrix_36_2 = 252'h9fc0059b29d98d4a1e898b1e84186ab754803dfd0e5ab54a92f006eb566456f;
  assign mdsMatrix_36_3 = 255'h700f4b271a6f81b713d6daf8b04b451fcd1dd8fa46a9602046ff7b18e0ce612c;
  assign mdsMatrix_36_4 = 255'h5bf3f52ac444f2cdf586c0e4bd1451a94cf8fea43101fc76c3fd90a5b215d016;
  assign mdsMatrix_36_5 = 252'hf31535f47129cbda4d2a2dd7cb59b38d8f24e7a81815b8f2c94ad1125b83209;
  assign mdsMatrix_36_6 = 254'h3c8188588cb3af2584639519c5866c9554e44d49c73fa6c81b0d92c6f40a99b8;
  assign mdsMatrix_36_7 = 253'h1395f154b79cbbeda47f11026ce0c0a4a12342985b328c5e0ab32d069ed7ca9c;
  assign mdsMatrix_36_8 = 253'h1dc602c49de6adabdb75e35239450448293c04f5cc495e801f9e80c663f18d6a;
  assign mdsMatrix_36_9 = 255'h42972d6c0ec56869e0573ee5d572b489a9c03f90f91f038ad4a54038ca935857;
  assign mdsMatrix_36_10 = 255'h582869ef815e40c2438f35de4a0fbfcfab532c661a937f14458d2ed1673ab900;
  assign mdsMatrix_36_11 = 254'h2c222391f8e7121d54bc9574525c07968ca90e7a0936b23acbff32c23c142d12;
  assign mdsMatrix_37_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_37_1 = 254'h3cf89c834f18d9555717e2130be3d5760d0fad89e3940ca6f25ea44c7902177d;
  assign mdsMatrix_37_2 = 255'h4947ed78be97e5b4c66f21d12181cab36a36453331970522e9ef78032ca14bf0;
  assign mdsMatrix_37_3 = 255'h44ec9ebc9ca617f1e111eb80d6d4db012b356908ed21131b5ea809fe53a745d8;
  assign mdsMatrix_37_4 = 254'h2ad05b66f92a437975fc1a5272b3b3cf956cde3cee9d4165349b217c3fc1f219;
  assign mdsMatrix_37_5 = 253'h1398f069acb9a7819e5c9f7a5806293b8e527e0090d944b644b1472998dc0edd;
  assign mdsMatrix_37_6 = 252'hd632b94dfea49ffb23f9c876012e6a8093b180eef997ca9a965200c4d4e2ee1;
  assign mdsMatrix_37_7 = 255'h663f055a034af952a022e725f21368dab8adbeeb9d25d285cecd064f526d8f5c;
  assign mdsMatrix_37_8 = 255'h72d1d6c8eb457cf339c1915041439d8c9e94a5012c0847cab3dbc4edd73de2b9;
  assign mdsMatrix_37_9 = 255'h4dee633e329bfde509af13a867e227d3b22ad37e72a1c3b062fc548401bc6509;
  assign mdsMatrix_37_10 = 250'h3ae2461a34659e0aece3ad7c7cdfce4243f986c1f049173b98887fce04443f7;
  assign mdsMatrix_37_11 = 251'h5dcb0413f6142205448f3e963bc09441de9a40828e9aaeed3e7b1ae58a26a9f;
  assign mdsMatrix_38_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_38_1 = 255'h62cabaaeba343fe2fc0676844038ad92fa523e5a8ce2fb88da39f481b626b18a;
  assign mdsMatrix_38_2 = 255'h618533f778f887951941a400241bb091b12b50e1f3056006cfa83b0c7938e37c;
  assign mdsMatrix_38_3 = 254'h30012ca0299b8a2740061d50c45d8b7fd902a604c51f457a5bf6400e631fa5f1;
  assign mdsMatrix_38_4 = 255'h527e53c960012b08bd1993efd40c5907733faafdc7c2032c140250a180bd7827;
  assign mdsMatrix_38_5 = 254'h3c909783c5f4491031b4c7de702df7c249ea37312465adfb2d10388836210d8a;
  assign mdsMatrix_38_6 = 253'h18998260a03c4afc303c15aa9f673b359399982dd44b4bc96ac0db1ebd7c8394;
  assign mdsMatrix_38_7 = 255'h6fd85eae9b9a23289f91a2b707040845ada7e5d0dd81dddc1ea09e25822c2728;
  assign mdsMatrix_38_8 = 254'h3c16034dd59b423d06dd3c59999fc6fbe780feedcad57c5bacb34553dd399855;
  assign mdsMatrix_38_9 = 255'h71647a58e128e9bd66dd680f540aec4988a5b133aecf1baa8a16be00a3d9e64f;
  assign mdsMatrix_38_10 = 255'h62df79f9c3cf566c9088d22c396fef2960f8adbfa80f2016556cf4b84cdab14f;
  assign mdsMatrix_38_11 = 254'h25746e20f23337419c0ac8f8c50084e248874a21ed8b57b13bd4f93977787545;
  assign mdsMatrix_39_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_39_1 = 255'h4e139de63123d5bdc985180adadfc5ec037554eb979f447f2bc7ef0815e56747;
  assign mdsMatrix_39_2 = 254'h313515a77ab8e3efd398f45a3c8d43d1905ee6c17bda4dc45de50cd8b4598100;
  assign mdsMatrix_39_3 = 252'h97d254f285220245e5d8647824d0728706b132f7a4e39dd614f79a350c67d17;
  assign mdsMatrix_39_4 = 252'hd02b90c15fe142e561b9f6d61ae98222a432a172f9b909b44969f7f6bcb927c;
  assign mdsMatrix_39_5 = 255'h50b764bdd6c2c1ffa0934d73e436a5595f57951f12bd762391b0f6169204a81c;
  assign mdsMatrix_39_6 = 255'h5d669b5ce88aa2c303b5de6dcfab677a6cfac69a4069e1a7bd27b0d2fdfbb273;
  assign mdsMatrix_39_7 = 255'h585a80611e31935fe825f0c51c154cd58181fbdfd116d46385500f89517352e1;
  assign mdsMatrix_39_8 = 249'h10192683c5adbb0b0d6b245eff94afe7786fee31b5dffbbf8ba26930714d389;
  assign mdsMatrix_39_9 = 254'h26a7a8eed0d286a0bce7cda93affc0972c94875468b5452278c608c139ff793f;
  assign mdsMatrix_39_10 = 252'h8cbae7580dbc7083cdd379c07e1e2d286113c100b73385e6b39e789ef927156;
  assign mdsMatrix_39_11 = 247'h7ced490ca0f7334d9b5accaa0ec5f833c769abe94efbfd9b5bcfe1c0b27233;
  assign mdsMatrix_40_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_40_1 = 255'h46717114d71919ac12007999e5bf0b279da63dcf82204f0c5b1fa603a47dcd35;
  assign mdsMatrix_40_2 = 254'h3ecf053cc0b2dd4fc09bbefef4673d64741e36d235d36d9050e09eeb728c83f4;
  assign mdsMatrix_40_3 = 254'h294d4bbcf810a7863c17ebc5ea18b586ce6e85ae91ddb7315ea9ec936ce3dfbb;
  assign mdsMatrix_40_4 = 253'h1a1b3e063047d31569079c598eea8f17205af26527207acbd1f110b8859b4b9b;
  assign mdsMatrix_40_5 = 252'heab89746f38bed2159f42ce93038a40a86cb8fa1ac0c44627fe944d84c72201;
  assign mdsMatrix_40_6 = 252'ha9d848fa780385c3ecd604b1574514972a571bdbe0d49eb6d49197a8bcd6f4b;
  assign mdsMatrix_40_7 = 254'h21b2bc8802a6494cac54217a7706dca9aff78e244ecfe561b13adc6690b30b63;
  assign mdsMatrix_40_8 = 253'h1631502c7b587abd61d36bd2f090b855b742372ff60047d46ab7ed1cee6aa92d;
  assign mdsMatrix_40_9 = 253'h1134d79d68c3cd4b55df2e40a20b7ba95c6ab8af43977f5e99245f436bfcf661;
  assign mdsMatrix_40_10 = 255'h40fea70f87ca24791177159c42348ede4924974f66cb39d756e7c2eabc6cbc87;
  assign mdsMatrix_40_11 = 253'h1d890c9b4a3901f44983d44c60f276dd59cbd39493b91a675508e48cea810c7a;
  assign mdsMatrix_41_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_41_1 = 254'h2ce01489c73b3ae8938b6aea0e284e91fd997b3542afdf2560edb29165ce851f;
  assign mdsMatrix_41_2 = 255'h596b8d4e79c75e9eb8fb20fee72c23c2ffca2df6c759fa85d90b8f8fcafcfb95;
  assign mdsMatrix_41_3 = 255'h538d722a6c94857e3acd6dd57e6c3394ad0899632837c042ab90321f6f815d29;
  assign mdsMatrix_41_4 = 254'h2618e5ba04e10ffff943fb7dc5c05618b719f579b56a0e69d871b2cea12e4a57;
  assign mdsMatrix_41_5 = 254'h26263a2cd724a5b2c7f3e44b7aaf34d4a4ab9250047488fca271dfa7f8483505;
  assign mdsMatrix_41_6 = 255'h4192ee56c1ca8c1f0be4cdf6afdff58b52b78a95b69f9b25638b9de1fc5a6fc4;
  assign mdsMatrix_41_7 = 254'h3edfdb7e62b945f313ddff5c28b655684ac5dd096500b04067239985a5a703f3;
  assign mdsMatrix_41_8 = 255'h6a0676d0f24a9f151d434e74f57eeb542499cbe157b9d06e50506593818c2a40;
  assign mdsMatrix_41_9 = 253'h1ddc4bf4d05ebf148f3372b2f2aedd69eff1cd0110ed4274ff797489001a0fcb;
  assign mdsMatrix_41_10 = 255'h4473da48be976346ae85660bb7978160937a03270ee602026dabe72366f93ad6;
  assign mdsMatrix_41_11 = 255'h694f846088426c0e1868e7d2b21d1333d0a5ff40ad8e59a146aa87102af75ea9;
  assign mdsMatrix_42_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_42_1 = 254'h2b72e2145926db5a6e4d7df2ae2c792fde54155959f6d1ee643f33d3df0059b9;
  assign mdsMatrix_42_2 = 254'h2d27c05fcde0d0e6c7ddbc4393c20e56456799105d33994f399ab6d7b6e91d5a;
  assign mdsMatrix_42_3 = 253'h1e35e5e37b6c388145d29c50cdd1f9dbf0611a7537edcd2d876f8efea1508740;
  assign mdsMatrix_42_4 = 255'h4caffd959d8fc20ed8c8d0b59ef7102efaf087caf85e8dff3fb6fe35213a0186;
  assign mdsMatrix_42_5 = 255'h49d71b6f4832e61148ae0ec08131f89e71733eb6a82d0e2bffcb32146c44f76e;
  assign mdsMatrix_42_6 = 251'h49d242697e747de361f3149caa3e4f1cd9686d9ea2e9007ebf09cd39b0c7a70;
  assign mdsMatrix_42_7 = 255'h6704d31ac67651fb59d63eade7300a383ce8001ae6b0f166d91b0f8221bdf56d;
  assign mdsMatrix_42_8 = 254'h35c8c03cb3f9637e0cf5b2447168cd4605739b7216532fc7b3eea63270244832;
  assign mdsMatrix_42_9 = 255'h44be45cbf3202effd72028b748307276441f08e1930be3908ab1fb93702f1363;
  assign mdsMatrix_42_10 = 253'h1de618ce92f1242b28b7f3ae6b8995ee2179c3220625886415ca4184af8f5d2e;
  assign mdsMatrix_42_11 = 255'h487933e61311337d318bf60907bb9dcbb3849102b283eba14e7dfc022ad15d93;
  assign mdsMatrix_43_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_43_1 = 255'h4968288cbdd1f065ec2596213415424693db64603d14d1df3f506bdce31880c6;
  assign mdsMatrix_43_2 = 255'h545c6a05a18d3d2e22b7cd10622843729125922a55db4a796f4ba63a450eb260;
  assign mdsMatrix_43_3 = 255'h648ffeda5c0ad9b9df2c8897bf81a61a1d3f68e6d97467c02760cc5ebcf69755;
  assign mdsMatrix_43_4 = 255'h71bda0a88930b276b2d09b30a25e17b9b16dc74f4ca4b826fb83c98eed20367b;
  assign mdsMatrix_43_5 = 255'h459d2aca86c8a569d2a96016cf852d415e4e9e3742e2e0e266370cc67792066c;
  assign mdsMatrix_43_6 = 250'h2ce01e2cb4c221bd40b94df6c2678b00d5fede26c352441280816549e004c32;
  assign mdsMatrix_43_7 = 255'h421f3a93fcb4be32360fd0b98bc2ff4dd13219a810998d7894e8d7f0ad965e6b;
  assign mdsMatrix_43_8 = 254'h3d6c7db5beb5156edccd0af5b4f957d9a586c6ff5047185bdc50228b60f5c54e;
  assign mdsMatrix_43_9 = 249'h176d835eacda85bed8efa3f488914c506572eaee3c1ae9d8cc17fe99b0aa175;
  assign mdsMatrix_43_10 = 255'h5415e5a1d31b5a30b914f8aec47dec343ccff4f7d63b4aa2fcbb96ce97a8bd86;
  assign mdsMatrix_43_11 = 254'h37e11453e5a824ca4e196b00545c385d2200c65517a770ffd5ca87fdc748b384;
  assign mdsMatrix_44_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_44_1 = 253'h1da3fc87bcbe89ca3d3f6858fb438edb79975e19e9c54392058fc9695584b767;
  assign mdsMatrix_44_2 = 254'h22a339441c7745e6f90af2a3782725ad811ae3573baa516b92d10768e45a480b;
  assign mdsMatrix_44_3 = 255'h71933b0c8a2926f8a16afede0a49ce49e96ddaa9e4e3fe7cfd22341f57c80111;
  assign mdsMatrix_44_4 = 254'h20ec1d5c315c3f6993798c3b9e44321adb7325ad4e280e9d119971cdd9da7751;
  assign mdsMatrix_44_5 = 255'h55f8d52706c89b5f9724b0963d53628456159eeb64a5f99535aa1bbe16e336bb;
  assign mdsMatrix_44_6 = 253'h1d776a6eb00009a8cef828652892ee0e52d4b6131aaf713acc8411bf1ad6d7d6;
  assign mdsMatrix_44_7 = 255'h7300f4fb94ee38f55ef8b07c4b8278caa2dce157e35dbc42e4e4616054760715;
  assign mdsMatrix_44_8 = 252'hd9e0955d6171d218ef605d8749affa7dd9c4af50b903b0b5460cb0a4290d147;
  assign mdsMatrix_44_9 = 254'h27ad4dd48a0fed127a3002a27fdba6dfe31e9aadb1a8df61ec4d69e89b1ed788;
  assign mdsMatrix_44_10 = 252'hb8e71eeee0cb8936e095d7eb275f3195f368b29acd1be86f6d3a601d7801fa6;
  assign mdsMatrix_44_11 = 255'h66de7583724fc06d4ca0b3566b33d95672566331b15d40907e63ef49975faeec;
  assign mdsMatrix_45_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_45_1 = 253'h10aec7e6a4c92cd843bd801f5e6559a48500fb3c06df995f94db0cc7b81e03d3;
  assign mdsMatrix_45_2 = 253'h1e33e532ecc728ecf53325198d7107325f448d41b14c8ce79d07b1d4e05e2635;
  assign mdsMatrix_45_3 = 255'h73457523cbfcf5dca4e3da5be11c9849e81637dec3accd25d42f81d189a2bffc;
  assign mdsMatrix_45_4 = 253'h177d7d4a84fe5b756f6bb4a11ceaa88fd6caf1c583f831978ece193fdecdb3d5;
  assign mdsMatrix_45_5 = 251'h4140dcaae13858b42c47b8ae71e84a61a009b965b0c4fcd0528dcb94781960b;
  assign mdsMatrix_45_6 = 255'h44eed32558b25b1a4ad2ed1c1a7f47bbebd4ae59e2e692e6c5c4f30b55a60e8b;
  assign mdsMatrix_45_7 = 254'h31aeac4c966182e1d525865b95aa6821d8e5a7ae5ff2ef51a7f7f9fb92a8c642;
  assign mdsMatrix_45_8 = 255'h63f776911b39c9ecc6ec8630ac87935c2069e8b53d881e0142535097fd89d0e6;
  assign mdsMatrix_45_9 = 253'h1205d3553995634781cdbbce7c321d06a3016520efe882abdffab81446f91d09;
  assign mdsMatrix_45_10 = 255'h63846452786d2398de7f065c29d652fce7576412261f89e19945d2eebdb21972;
  assign mdsMatrix_45_11 = 255'h57bfe3bf3bcbdd62aa997609c6de85ff5f035ad7a0f30c4c0ddd5f33eee61179;
  assign mdsMatrix_46_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_46_1 = 252'hea57cbc152761ac519d5db2a320fcc9beeeb85ea7e7aa79dfdd80880a2df4c1;
  assign mdsMatrix_46_2 = 255'h58305cd24117bba0856df0e9d857d4fec814fd95f3992e00c5440bb675c09aa3;
  assign mdsMatrix_46_3 = 254'h37d2e6bc314d25fde499b25917784323061c35610e051fa93b89bec0147970ba;
  assign mdsMatrix_46_4 = 255'h550278ad6a72da480050d1c3516e89686fd29316c0f156dae6031ec4aab83839;
  assign mdsMatrix_46_5 = 255'h5ec79dda32f4e9e5b451abcbb3891b58b4eb3e8313f7e35c20f0bd7b47085d72;
  assign mdsMatrix_46_6 = 253'h1100c47f421672b78481151464ffdf4c20c26f824fc55fb44623a3a8eb65ee3e;
  assign mdsMatrix_46_7 = 253'h1c1496a842ed55c67c70ef2c765809ebb845b24a1d70b4ae512322274fe4b524;
  assign mdsMatrix_46_8 = 253'h163d31b6307a8516c80f59b0b8e4c676f04579403cf10f1509a4f331b879c801;
  assign mdsMatrix_46_9 = 255'h58c9bb4a436b8d27fa269a246a69bd276d5a25b3ecd8214e087147d218268a8e;
  assign mdsMatrix_46_10 = 255'h517b46748017a07f910d45b3488aa9c5b4354d9a63f7ef0c1e0f9c4c4f094b66;
  assign mdsMatrix_46_11 = 255'h49dfef83c146c0cee7359b8b5992e63b7ef1ea8aaf0a13efde8ffb7cd8db993d;
  assign mdsMatrix_47_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_47_1 = 254'h2adf512069e204eb38d0b1a1d122989f9bd2468180e78357d0b1473ff4b62bd9;
  assign mdsMatrix_47_2 = 253'h1eecc9e53528ae97138b4620aa927598fb4dc83be0e0a50dbe22c174cc7fbd8a;
  assign mdsMatrix_47_3 = 255'h43ed70f9800e1b231f6c3eafb6b71f9236974e5b96583cf8b08a8f9e4aff275f;
  assign mdsMatrix_47_4 = 255'h51466f94805ecc2d8f52ecfe7f72aa0caafd03789503e05640bbcd2e953317ed;
  assign mdsMatrix_47_5 = 254'h3aea683becad8a0f514e965faade1ea86148ca945ece6016b99e01696b1f2aeb;
  assign mdsMatrix_47_6 = 253'h103154683ce17fbed07127e8f8e4d597af3abf471217d8a6edcef55e0cc79484;
  assign mdsMatrix_47_7 = 255'h4ad091e6dbd55addb652d696c4d4ce6d21dfd983d5c2ae4daf5ac393fd744197;
  assign mdsMatrix_47_8 = 255'h4cf8a6bf2b7a20e34008d3deb56b0f1698f89919c73594abd235216b3de914ca;
  assign mdsMatrix_47_9 = 249'h152247f6c7825506d9206e349e3d92a739fc24452ce6aa13986e4a14fc1c345;
  assign mdsMatrix_47_10 = 255'h46f393134e136eb6c1ec1ee6e3b0266c5ec3fbe48ff928721515f1a6571d4e40;
  assign mdsMatrix_47_11 = 255'h4a949f8a204f9be6846f27322dc2ce299d2bb4a9b8d94f49963612447905e2bc;
  assign mdsMatrix_48_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_48_1 = 255'h5b242330db8a26135035edd54544e0de72a0b616bf92e8413b613810b972da24;
  assign mdsMatrix_48_2 = 255'h5e910f10a02d369e8775f302bc0c98e5d604cc22ae4da1d96d9046c1112ef35b;
  assign mdsMatrix_48_3 = 253'h1d61af76e9e45c1cb895ee03d79756f92bb603a13a636d9d9be3b186e5c3ee2e;
  assign mdsMatrix_48_4 = 255'h66c2785311b2e990073013d7e99d6a6dd58bf0303c52f9391ab229cafe6284a2;
  assign mdsMatrix_48_5 = 255'h4dc39d9729428bde63739efaeb5744069b28a4db82ecca723bf18c0b08d611ff;
  assign mdsMatrix_48_6 = 252'hbe8f2eab4f4de00c3abc04292c6df00b093115b47a79888d39b9007b414d163;
  assign mdsMatrix_48_7 = 255'h5f595b093b4c837567f989bba2ba6dc5b3e4460e818d25982a82397008679df6;
  assign mdsMatrix_48_8 = 255'h4470d71d7b516402241d2715651b8c45c02d42ac15db9308c35929594e6dc1c2;
  assign mdsMatrix_48_9 = 255'h6754bf508a33394afcfff5b75c8cd989b82d9bff2e076b059e1a4cdae8d08311;
  assign mdsMatrix_48_10 = 255'h50f0c44bba71255401f8f0d0d2b24a1f47c2691040c5c42698ea8ee73c5a6177;
  assign mdsMatrix_48_11 = 255'h6f871409d3295515a85ce926ee63b99ff851e5b08b064fb6d09ebe3aa06f93ce;
  assign mdsMatrix_49_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_49_1 = 251'h44274e9a774cf50d03fab1096dcc6cf5542b3dc43d0df94d1eb75df1914d555;
  assign mdsMatrix_49_2 = 255'h5a5d6ffca25cea48e48885faa25c198f6971305ce5ba74d204833c15ec0e0f45;
  assign mdsMatrix_49_3 = 255'h43c26f0f894fc5f1699fb8e29e16a4524c3bc330a674dac4e8982be4aea4fe4c;
  assign mdsMatrix_49_4 = 255'h4c0272e315f9025cb51c0a4d1a71a42a8455f434408b59263437ccd25506e9e7;
  assign mdsMatrix_49_5 = 254'h365e7c01f60d8bb4a183fb1f9d867c49910ff19a18acc140b943d1228fef3508;
  assign mdsMatrix_49_6 = 255'h6cd30a9c6346586c01f7834728d76b9aa2a736157f95ea8efe1c6ecf897d076e;
  assign mdsMatrix_49_7 = 251'h459090c5bc3db616d6a634fcb76008a692874e54894c085998146f966bcadae;
  assign mdsMatrix_49_8 = 254'h204cf5510245bbb15792f1ed5609a800429f1f9b08767922e55a26a924e65f81;
  assign mdsMatrix_49_9 = 255'h46ccd8a16b6a264b1fe44e860c76fb117b91332e495a0e349662aad11c569c1a;
  assign mdsMatrix_49_10 = 252'he44b5a8ae53295d211e7b61c09ac90fdd368b9f7795830d29963f7a474bdf4c;
  assign mdsMatrix_49_11 = 255'h68307048c2bd7f528a4558a302fb92aa4e8be2bed68d162ef0ab5853c3bddf86;
  assign mdsMatrix_50_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_50_1 = 255'h6973f64f6e38c8da454ea4a39d284e6d63846ec9225ee536899d1d443d336c73;
  assign mdsMatrix_50_2 = 254'h2ee730b2f04ff130d0e868d4d001d40c55ce44b7f31b15a86f51a67d32c14a14;
  assign mdsMatrix_50_3 = 255'h6d90135f413c927698f9a784bf6030f67d8147214a582983d066c49d1273c9b5;
  assign mdsMatrix_50_4 = 255'h614da2f5fcba16ce67f92e074ad78c4403c8e3b14760b98783874af229a52cef;
  assign mdsMatrix_50_5 = 252'h992fd477855368478aea6d6897d0384ea9843335f8e0075357222ff59852536;
  assign mdsMatrix_50_6 = 255'h650816f12d21a4205cd5c34316fcada3dda715eb4b2a474951633b0d07c6fad3;
  assign mdsMatrix_50_7 = 255'h58862a1622ef2ccea93272b2c19b50b0e54fd3b33581614d8a2decf163b3aa35;
  assign mdsMatrix_50_8 = 253'h1a9c4b5b577c628cb5c9fa455440de807ef3e7c9ec535dceab8c8a5d85832155;
  assign mdsMatrix_50_9 = 253'h1f34ef34c07d73686a2009e063f55ed76ddeef6b7406e2ae75de4a7c1fcb5602;
  assign mdsMatrix_50_10 = 255'h56bf547ce770a9cd3470b1db85ce2c6a8e09f26ed424ab76d0d3b054322c3bd3;
  assign mdsMatrix_50_11 = 255'h4506dd7f143354b98529b9c29d7b31c0372564b64607113c10825c383c7ae8b1;
  assign mdsMatrix_51_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_51_1 = 255'h73ed2e22d11c8a677851d9973ad8c2fdbf698b04c368b2fbedc60bd3e94b3ff1;
  assign mdsMatrix_51_2 = 255'h49315c95b84f07b875eb485339bd77905f7c0203137bcfa63cf7a1277dfe32d2;
  assign mdsMatrix_51_3 = 254'h2ded93b8de954a3b6bc2fe7cf16c60c1958dd684262dd7776d866f33d8f25a0e;
  assign mdsMatrix_51_4 = 255'h4a9cf2e16fd1e69a73301f25556cfa6c41acbd379bb393f8b4332ba7deec3f6c;
  assign mdsMatrix_51_5 = 253'h1c8befbe4df735ddbe89cddfda4396de69ed252d38d2a47c16cc47df126ebef1;
  assign mdsMatrix_51_6 = 255'h6237ab62b69afb80f97f094c51d5785b4a15ecd716cb456e806585722c837e70;
  assign mdsMatrix_51_7 = 255'h50dc99edf95e3b77ecc06e026ee2855b0645b4ab2d98abbaf4ea5cbd9fa7f716;
  assign mdsMatrix_51_8 = 254'h334a0b48d283a169f0696d30ad380dece7240a12bb06aeb12fd4399111879cec;
  assign mdsMatrix_51_9 = 255'h5ce8ec1c64095eb997caa42c3672f73fe3e957db9f15f233be6eb7e72441489a;
  assign mdsMatrix_51_10 = 254'h32e612bd13bab65915c0dccc0bf3c019012df08bc6c11a5f3ddea5c8c5a0a0a8;
  assign mdsMatrix_51_11 = 255'h438cd76de72011a3bf29664cb540d8e3cccd14922b8ee7f9ee5829ac7bad2a8e;
  assign mdsMatrix_52_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_52_1 = 255'h5adfafc3fb68647139b0ad8a9777770833439440b899cf1f4fff5a96ebef7cc6;
  assign mdsMatrix_52_2 = 254'h2b1acb3d0d9af933a7200cf7906a44e5c51ad25b0cbec53677b6f431f5616f2d;
  assign mdsMatrix_52_3 = 254'h21eb58fc2a59add1a5129fd838af1b896b6a06f1c9759531fcc30329749b2e9d;
  assign mdsMatrix_52_4 = 253'h11b32338626d331089319fefd0d683f99df88a2e39462742196ede27e402dcd8;
  assign mdsMatrix_52_5 = 254'h3a30eba49b49836ec96590813dc6be4119d482d872d3fb561a1bccfbc4e6e58b;
  assign mdsMatrix_52_6 = 255'h6d2129b10a4e17e104184ce5d8aed76fdc6db0e9356813e3dfeaf67e2006cb29;
  assign mdsMatrix_52_7 = 255'h6bf71b846147d9dfb573448c23aef981cfdc94b1cc73cf07402dbdb5cb547272;
  assign mdsMatrix_52_8 = 254'h224f170c4bca3d313f95ceaea0a72ea3174b71a8d4c2605e9bb0a2415dcb72cd;
  assign mdsMatrix_52_9 = 255'h4040cfc89ff924042e8accc7d8db475c9cda9813779d30c8a954a6fa631cf751;
  assign mdsMatrix_52_10 = 244'h8688d6025290b13b219add3959e0baaa7ade196e04d48895be5c528a99db2;
  assign mdsMatrix_52_11 = 255'h5340e409534e45d620a573f0994a29a3e3c90bc718620a18149541a63a87f116;
  assign mdsMatrix_53_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_53_1 = 255'h4057301ec03ed106cb5b71d5b9028e30a36ad647ef9302481def551ebef4cfbc;
  assign mdsMatrix_53_2 = 253'h1d179f007ae0ebbc08ec155582028dd2197e523890d12d559fce54f6f0708a31;
  assign mdsMatrix_53_3 = 255'h4e43d30d13a8798429e1bfef2f7fb8ac17bd490aecef8ea78e175553a7c81934;
  assign mdsMatrix_53_4 = 251'h63cc0e8d0e8b115a0e0cdd4c43bb65ad0e5af9e27f5ed6c69df86d9cdf334b4;
  assign mdsMatrix_53_5 = 254'h2194b1c417ed54f1e395c91ecac0394f3a532405ebc44fe067c52314466d7bf1;
  assign mdsMatrix_53_6 = 254'h2e0d93a324bdffcdd1be5a2fc1d66bc33fbbdc3daa8b2b709588ee1180e77278;
  assign mdsMatrix_53_7 = 249'h11ef27c5e234d48416374236df7106a59af3d3c5c092feb3e38ea74053c4270;
  assign mdsMatrix_53_8 = 253'h17c4ed37b9a2f0417e652967bd7b08f95faae414c09c2094c6d6dcf0b70aa25b;
  assign mdsMatrix_53_9 = 252'hb2adc28c854f48136f9882ba27bf109d65fc2532b1b5f14a9f689df665a5ea2;
  assign mdsMatrix_53_10 = 255'h70c651b309b764fc0f829c11922b83a54ccb64b84b13889e083bcc71776a406d;
  assign mdsMatrix_53_11 = 255'h487a1b61436cd5b9b2a0396ccf7284c79e17db3ff6b438763907327378de4ef2;
  assign mdsMatrix_54_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_54_1 = 254'h3812db2ffe6e4fb7dcca194bbe31c59b37006b76696fec1556b4fd6c0d950cdd;
  assign mdsMatrix_54_2 = 255'h4e294b50951adf3c3f919db6ccbfe436db4e1a1d384750487a5f5789eb622048;
  assign mdsMatrix_54_3 = 254'h38022e7949e9c5cbf5dde8388b2216c502289664ba69379bd25474717182eb23;
  assign mdsMatrix_54_4 = 252'hf7194e41da09f76c3ab74f23281fa71bf26079e2a214d2e62321ec1109e2821;
  assign mdsMatrix_54_5 = 254'h3bb700ca2e04e83b0443cc82f1e57df85da40468528064626f88b907544efd3d;
  assign mdsMatrix_54_6 = 254'h2169e5bc0ca788d24052ebca303c085673dc756a1f3d4a54fc0c03029a5103db;
  assign mdsMatrix_54_7 = 255'h64a1a03a8ae2f0f040915293416184c3f7cde255e1a5c343eba0d713db0b1578;
  assign mdsMatrix_54_8 = 255'h4c9129ef609d9e7e5760d5209d3b4684d7ae8d559af3b4cdd1339744b50d0fb6;
  assign mdsMatrix_54_9 = 253'h1e90bf90d75e64482c2f1bf9be41788d68001d22998bfe9498b03af3b58cd583;
  assign mdsMatrix_54_10 = 255'h5f43291335ed3fa19685af1e7f814a9e7c15f2bdc836f7699ebe79b780b0edc1;
  assign mdsMatrix_54_11 = 254'h284ebda357391a381b19c72a0d7b78b0b6ad730698136b659f02a0c6eeb97fcd;
  assign mdsMatrix_55_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_55_1 = 254'h20ce49b5295b61e76cf82c506b0060d324deb20dbe5b8f96c4ec4ec4b7cb7cb8;
  assign mdsMatrix_55_2 = 255'h57fed3e9682e0e741a8f2c35abc1438878a35decd378e48be61e61e56eea21d6;
  assign mdsMatrix_55_3 = 254'h33f4687c8f33241b16de2e9e8dc0b292935bcfb2373607b8cdecdecd8c058d26;
  assign mdsMatrix_55_4 = 255'h4035f07319cd8c4db0eb4ef88d763b6a46b03acfc11c562936e36e3666a55945;
  assign mdsMatrix_55_5 = 255'h6510f90b93578087d2bb119f9c5a7692a0015902ac204f080756dbd354b2bf07;
  assign mdsMatrix_55_6 = 254'h2c2ef123dc3b7b06c53e643d056e98d0e8bf4cbe4e8aaa5d31c37a6086027b8d;
  assign mdsMatrix_55_7 = 254'h355646ee2b6b9b267a769661368415b2d8519c1552973da077a5a0b6b28337fc;
  assign mdsMatrix_55_8 = 254'h2c9eb19d62935f8f50cfbf87aabc4e8573f4acb6eccf1bb0f9350da8240b2d7a;
  assign mdsMatrix_55_9 = 252'h83b6bc7a43728fdd01676f049435226992cc31642ec04b8acc171ba4e177b0c;
  assign mdsMatrix_55_10 = 255'h421cbc273523c66f26807150aa14350c980de30d02d20a2fca0689431949e255;
  assign mdsMatrix_55_11 = 255'h4fcf2780f2571f771150f634c56a7e8a0c4bd03bd3d6c6ead0f4bd8abea91141;
  assign mdsMatrix_56_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_56_1 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_56_2 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_56_3 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_56_4 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_56_5 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_56_6 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_56_7 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_56_8 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_56_9 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_56_10 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_56_11 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign tempAddrVec_5 = io_addr_regNext_5;
  assign tempAddrVec_6 = io_addr_regNext_6;
  assign tempAddrVec_7 = io_addr_regNext_7;
  assign tempAddrVec_8 = io_addr_regNext_8;
  assign tempAddrVec_9 = io_addr_regNext_9;
  assign tempAddrVec_10 = io_addr_regNext_10;
  assign tempAddrVec_11 = io_addr_regNext_11;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  assign io_data_5 = _zz_mdsMem_5_port0;
  assign io_data_6 = _zz_mdsMem_6_port0;
  assign io_data_7 = _zz_mdsMem_7_port0;
  assign io_data_8 = _zz_mdsMem_8_port0;
  assign io_data_9 = _zz_mdsMem_9_port0;
  assign io_data_10 = _zz_mdsMem_10_port0;
  assign io_data_11 = _zz_mdsMem_11_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
    io_addr_regNext_5 <= io_addr;
    io_addr_regNext_6 <= io_addr;
    io_addr_regNext_7 <= io_addr;
    io_addr_regNext_8 <= io_addr;
    io_addr_regNext_9 <= io_addr;
    io_addr_regNext_10 <= io_addr;
    io_addr_regNext_11 <= io_addr;
  end


endmodule

module MatrixConstantMem_10 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  input      [5:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  reg        [254:0]  _zz_mdsMem_5_port0;
  reg        [254:0]  _zz_mdsMem_6_port0;
  reg        [254:0]  _zz_mdsMem_7_port0;
  reg        [254:0]  _zz_mdsMem_8_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire                _zz_mdsMem_5_port;
  wire                _zz_io_data_5;
  wire                _zz_mdsMem_6_port;
  wire                _zz_io_data_6;
  wire                _zz_mdsMem_7_port;
  wire                _zz_io_data_7;
  wire                _zz_mdsMem_8_port;
  wire                _zz_io_data_8;
  wire       [254:0]  mdsMatrix_0_0;
  wire       [251:0]  mdsMatrix_0_1;
  wire       [253:0]  mdsMatrix_0_2;
  wire       [252:0]  mdsMatrix_0_3;
  wire       [253:0]  mdsMatrix_0_4;
  wire       [253:0]  mdsMatrix_0_5;
  wire       [252:0]  mdsMatrix_0_6;
  wire       [254:0]  mdsMatrix_0_7;
  wire       [251:0]  mdsMatrix_0_8;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [254:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [254:0]  mdsMatrix_1_3;
  wire       [254:0]  mdsMatrix_1_4;
  wire       [250:0]  mdsMatrix_1_5;
  wire       [254:0]  mdsMatrix_1_6;
  wire       [252:0]  mdsMatrix_1_7;
  wire       [252:0]  mdsMatrix_1_8;
  wire       [254:0]  mdsMatrix_2_0;
  wire       [253:0]  mdsMatrix_2_1;
  wire       [252:0]  mdsMatrix_2_2;
  wire       [254:0]  mdsMatrix_2_3;
  wire       [253:0]  mdsMatrix_2_4;
  wire       [253:0]  mdsMatrix_2_5;
  wire       [254:0]  mdsMatrix_2_6;
  wire       [253:0]  mdsMatrix_2_7;
  wire       [254:0]  mdsMatrix_2_8;
  wire       [254:0]  mdsMatrix_3_0;
  wire       [254:0]  mdsMatrix_3_1;
  wire       [253:0]  mdsMatrix_3_2;
  wire       [254:0]  mdsMatrix_3_3;
  wire       [252:0]  mdsMatrix_3_4;
  wire       [254:0]  mdsMatrix_3_5;
  wire       [253:0]  mdsMatrix_3_6;
  wire       [253:0]  mdsMatrix_3_7;
  wire       [254:0]  mdsMatrix_3_8;
  wire       [254:0]  mdsMatrix_4_0;
  wire       [254:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [254:0]  mdsMatrix_4_3;
  wire       [254:0]  mdsMatrix_4_4;
  wire       [252:0]  mdsMatrix_4_5;
  wire       [252:0]  mdsMatrix_4_6;
  wire       [250:0]  mdsMatrix_4_7;
  wire       [254:0]  mdsMatrix_4_8;
  wire       [254:0]  mdsMatrix_5_0;
  wire       [252:0]  mdsMatrix_5_1;
  wire       [254:0]  mdsMatrix_5_2;
  wire       [254:0]  mdsMatrix_5_3;
  wire       [254:0]  mdsMatrix_5_4;
  wire       [254:0]  mdsMatrix_5_5;
  wire       [254:0]  mdsMatrix_5_6;
  wire       [250:0]  mdsMatrix_5_7;
  wire       [254:0]  mdsMatrix_5_8;
  wire       [254:0]  mdsMatrix_6_0;
  wire       [253:0]  mdsMatrix_6_1;
  wire       [253:0]  mdsMatrix_6_2;
  wire       [254:0]  mdsMatrix_6_3;
  wire       [254:0]  mdsMatrix_6_4;
  wire       [252:0]  mdsMatrix_6_5;
  wire       [247:0]  mdsMatrix_6_6;
  wire       [254:0]  mdsMatrix_6_7;
  wire       [254:0]  mdsMatrix_6_8;
  wire       [254:0]  mdsMatrix_7_0;
  wire       [252:0]  mdsMatrix_7_1;
  wire       [254:0]  mdsMatrix_7_2;
  wire       [252:0]  mdsMatrix_7_3;
  wire       [251:0]  mdsMatrix_7_4;
  wire       [253:0]  mdsMatrix_7_5;
  wire       [253:0]  mdsMatrix_7_6;
  wire       [251:0]  mdsMatrix_7_7;
  wire       [252:0]  mdsMatrix_7_8;
  wire       [254:0]  mdsMatrix_8_0;
  wire       [254:0]  mdsMatrix_8_1;
  wire       [254:0]  mdsMatrix_8_2;
  wire       [253:0]  mdsMatrix_8_3;
  wire       [252:0]  mdsMatrix_8_4;
  wire       [253:0]  mdsMatrix_8_5;
  wire       [254:0]  mdsMatrix_8_6;
  wire       [252:0]  mdsMatrix_8_7;
  wire       [253:0]  mdsMatrix_8_8;
  wire       [254:0]  mdsMatrix_9_0;
  wire       [251:0]  mdsMatrix_9_1;
  wire       [253:0]  mdsMatrix_9_2;
  wire       [254:0]  mdsMatrix_9_3;
  wire       [254:0]  mdsMatrix_9_4;
  wire       [253:0]  mdsMatrix_9_5;
  wire       [254:0]  mdsMatrix_9_6;
  wire       [254:0]  mdsMatrix_9_7;
  wire       [253:0]  mdsMatrix_9_8;
  wire       [254:0]  mdsMatrix_10_0;
  wire       [249:0]  mdsMatrix_10_1;
  wire       [254:0]  mdsMatrix_10_2;
  wire       [253:0]  mdsMatrix_10_3;
  wire       [249:0]  mdsMatrix_10_4;
  wire       [252:0]  mdsMatrix_10_5;
  wire       [254:0]  mdsMatrix_10_6;
  wire       [252:0]  mdsMatrix_10_7;
  wire       [252:0]  mdsMatrix_10_8;
  wire       [254:0]  mdsMatrix_11_0;
  wire       [251:0]  mdsMatrix_11_1;
  wire       [251:0]  mdsMatrix_11_2;
  wire       [251:0]  mdsMatrix_11_3;
  wire       [254:0]  mdsMatrix_11_4;
  wire       [254:0]  mdsMatrix_11_5;
  wire       [253:0]  mdsMatrix_11_6;
  wire       [253:0]  mdsMatrix_11_7;
  wire       [254:0]  mdsMatrix_11_8;
  wire       [254:0]  mdsMatrix_12_0;
  wire       [254:0]  mdsMatrix_12_1;
  wire       [252:0]  mdsMatrix_12_2;
  wire       [250:0]  mdsMatrix_12_3;
  wire       [252:0]  mdsMatrix_12_4;
  wire       [253:0]  mdsMatrix_12_5;
  wire       [254:0]  mdsMatrix_12_6;
  wire       [252:0]  mdsMatrix_12_7;
  wire       [254:0]  mdsMatrix_12_8;
  wire       [254:0]  mdsMatrix_13_0;
  wire       [252:0]  mdsMatrix_13_1;
  wire       [254:0]  mdsMatrix_13_2;
  wire       [249:0]  mdsMatrix_13_3;
  wire       [254:0]  mdsMatrix_13_4;
  wire       [254:0]  mdsMatrix_13_5;
  wire       [253:0]  mdsMatrix_13_6;
  wire       [251:0]  mdsMatrix_13_7;
  wire       [253:0]  mdsMatrix_13_8;
  wire       [254:0]  mdsMatrix_14_0;
  wire       [250:0]  mdsMatrix_14_1;
  wire       [252:0]  mdsMatrix_14_2;
  wire       [254:0]  mdsMatrix_14_3;
  wire       [253:0]  mdsMatrix_14_4;
  wire       [253:0]  mdsMatrix_14_5;
  wire       [250:0]  mdsMatrix_14_6;
  wire       [254:0]  mdsMatrix_14_7;
  wire       [254:0]  mdsMatrix_14_8;
  wire       [254:0]  mdsMatrix_15_0;
  wire       [254:0]  mdsMatrix_15_1;
  wire       [251:0]  mdsMatrix_15_2;
  wire       [254:0]  mdsMatrix_15_3;
  wire       [253:0]  mdsMatrix_15_4;
  wire       [252:0]  mdsMatrix_15_5;
  wire       [253:0]  mdsMatrix_15_6;
  wire       [254:0]  mdsMatrix_15_7;
  wire       [254:0]  mdsMatrix_15_8;
  wire       [254:0]  mdsMatrix_16_0;
  wire       [254:0]  mdsMatrix_16_1;
  wire       [254:0]  mdsMatrix_16_2;
  wire       [254:0]  mdsMatrix_16_3;
  wire       [253:0]  mdsMatrix_16_4;
  wire       [253:0]  mdsMatrix_16_5;
  wire       [254:0]  mdsMatrix_16_6;
  wire       [254:0]  mdsMatrix_16_7;
  wire       [253:0]  mdsMatrix_16_8;
  wire       [254:0]  mdsMatrix_17_0;
  wire       [253:0]  mdsMatrix_17_1;
  wire       [254:0]  mdsMatrix_17_2;
  wire       [252:0]  mdsMatrix_17_3;
  wire       [253:0]  mdsMatrix_17_4;
  wire       [253:0]  mdsMatrix_17_5;
  wire       [253:0]  mdsMatrix_17_6;
  wire       [251:0]  mdsMatrix_17_7;
  wire       [252:0]  mdsMatrix_17_8;
  wire       [254:0]  mdsMatrix_18_0;
  wire       [253:0]  mdsMatrix_18_1;
  wire       [250:0]  mdsMatrix_18_2;
  wire       [254:0]  mdsMatrix_18_3;
  wire       [250:0]  mdsMatrix_18_4;
  wire       [254:0]  mdsMatrix_18_5;
  wire       [254:0]  mdsMatrix_18_6;
  wire       [251:0]  mdsMatrix_18_7;
  wire       [254:0]  mdsMatrix_18_8;
  wire       [254:0]  mdsMatrix_19_0;
  wire       [248:0]  mdsMatrix_19_1;
  wire       [251:0]  mdsMatrix_19_2;
  wire       [251:0]  mdsMatrix_19_3;
  wire       [253:0]  mdsMatrix_19_4;
  wire       [254:0]  mdsMatrix_19_5;
  wire       [253:0]  mdsMatrix_19_6;
  wire       [254:0]  mdsMatrix_19_7;
  wire       [253:0]  mdsMatrix_19_8;
  wire       [254:0]  mdsMatrix_20_0;
  wire       [254:0]  mdsMatrix_20_1;
  wire       [254:0]  mdsMatrix_20_2;
  wire       [253:0]  mdsMatrix_20_3;
  wire       [254:0]  mdsMatrix_20_4;
  wire       [252:0]  mdsMatrix_20_5;
  wire       [254:0]  mdsMatrix_20_6;
  wire       [252:0]  mdsMatrix_20_7;
  wire       [253:0]  mdsMatrix_20_8;
  wire       [254:0]  mdsMatrix_21_0;
  wire       [254:0]  mdsMatrix_21_1;
  wire       [254:0]  mdsMatrix_21_2;
  wire       [254:0]  mdsMatrix_21_3;
  wire       [250:0]  mdsMatrix_21_4;
  wire       [252:0]  mdsMatrix_21_5;
  wire       [253:0]  mdsMatrix_21_6;
  wire       [254:0]  mdsMatrix_21_7;
  wire       [253:0]  mdsMatrix_21_8;
  wire       [254:0]  mdsMatrix_22_0;
  wire       [251:0]  mdsMatrix_22_1;
  wire       [253:0]  mdsMatrix_22_2;
  wire       [254:0]  mdsMatrix_22_3;
  wire       [254:0]  mdsMatrix_22_4;
  wire       [253:0]  mdsMatrix_22_5;
  wire       [254:0]  mdsMatrix_22_6;
  wire       [251:0]  mdsMatrix_22_7;
  wire       [253:0]  mdsMatrix_22_8;
  wire       [254:0]  mdsMatrix_23_0;
  wire       [252:0]  mdsMatrix_23_1;
  wire       [252:0]  mdsMatrix_23_2;
  wire       [253:0]  mdsMatrix_23_3;
  wire       [254:0]  mdsMatrix_23_4;
  wire       [253:0]  mdsMatrix_23_5;
  wire       [248:0]  mdsMatrix_23_6;
  wire       [254:0]  mdsMatrix_23_7;
  wire       [254:0]  mdsMatrix_23_8;
  wire       [254:0]  mdsMatrix_24_0;
  wire       [254:0]  mdsMatrix_24_1;
  wire       [252:0]  mdsMatrix_24_2;
  wire       [254:0]  mdsMatrix_24_3;
  wire       [252:0]  mdsMatrix_24_4;
  wire       [253:0]  mdsMatrix_24_5;
  wire       [254:0]  mdsMatrix_24_6;
  wire       [250:0]  mdsMatrix_24_7;
  wire       [254:0]  mdsMatrix_24_8;
  wire       [254:0]  mdsMatrix_25_0;
  wire       [253:0]  mdsMatrix_25_1;
  wire       [254:0]  mdsMatrix_25_2;
  wire       [253:0]  mdsMatrix_25_3;
  wire       [250:0]  mdsMatrix_25_4;
  wire       [254:0]  mdsMatrix_25_5;
  wire       [254:0]  mdsMatrix_25_6;
  wire       [248:0]  mdsMatrix_25_7;
  wire       [250:0]  mdsMatrix_25_8;
  wire       [254:0]  mdsMatrix_26_0;
  wire       [254:0]  mdsMatrix_26_1;
  wire       [254:0]  mdsMatrix_26_2;
  wire       [253:0]  mdsMatrix_26_3;
  wire       [254:0]  mdsMatrix_26_4;
  wire       [254:0]  mdsMatrix_26_5;
  wire       [249:0]  mdsMatrix_26_6;
  wire       [254:0]  mdsMatrix_26_7;
  wire       [253:0]  mdsMatrix_26_8;
  wire       [254:0]  mdsMatrix_27_0;
  wire       [254:0]  mdsMatrix_27_1;
  wire       [252:0]  mdsMatrix_27_2;
  wire       [253:0]  mdsMatrix_27_3;
  wire       [254:0]  mdsMatrix_27_4;
  wire       [252:0]  mdsMatrix_27_5;
  wire       [247:0]  mdsMatrix_27_6;
  wire       [254:0]  mdsMatrix_27_7;
  wire       [253:0]  mdsMatrix_27_8;
  wire       [254:0]  mdsMatrix_28_0;
  wire       [254:0]  mdsMatrix_28_1;
  wire       [251:0]  mdsMatrix_28_2;
  wire       [254:0]  mdsMatrix_28_3;
  wire       [250:0]  mdsMatrix_28_4;
  wire       [252:0]  mdsMatrix_28_5;
  wire       [254:0]  mdsMatrix_28_6;
  wire       [254:0]  mdsMatrix_28_7;
  wire       [254:0]  mdsMatrix_28_8;
  wire       [254:0]  mdsMatrix_29_0;
  wire       [254:0]  mdsMatrix_29_1;
  wire       [253:0]  mdsMatrix_29_2;
  wire       [249:0]  mdsMatrix_29_3;
  wire       [254:0]  mdsMatrix_29_4;
  wire       [254:0]  mdsMatrix_29_5;
  wire       [254:0]  mdsMatrix_29_6;
  wire       [254:0]  mdsMatrix_29_7;
  wire       [253:0]  mdsMatrix_29_8;
  wire       [254:0]  mdsMatrix_30_0;
  wire       [251:0]  mdsMatrix_30_1;
  wire       [250:0]  mdsMatrix_30_2;
  wire       [252:0]  mdsMatrix_30_3;
  wire       [254:0]  mdsMatrix_30_4;
  wire       [252:0]  mdsMatrix_30_5;
  wire       [254:0]  mdsMatrix_30_6;
  wire       [254:0]  mdsMatrix_30_7;
  wire       [251:0]  mdsMatrix_30_8;
  wire       [254:0]  mdsMatrix_31_0;
  wire       [254:0]  mdsMatrix_31_1;
  wire       [254:0]  mdsMatrix_31_2;
  wire       [251:0]  mdsMatrix_31_3;
  wire       [254:0]  mdsMatrix_31_4;
  wire       [253:0]  mdsMatrix_31_5;
  wire       [254:0]  mdsMatrix_31_6;
  wire       [253:0]  mdsMatrix_31_7;
  wire       [253:0]  mdsMatrix_31_8;
  wire       [254:0]  mdsMatrix_32_0;
  wire       [254:0]  mdsMatrix_32_1;
  wire       [254:0]  mdsMatrix_32_2;
  wire       [254:0]  mdsMatrix_32_3;
  wire       [248:0]  mdsMatrix_32_4;
  wire       [251:0]  mdsMatrix_32_5;
  wire       [254:0]  mdsMatrix_32_6;
  wire       [253:0]  mdsMatrix_32_7;
  wire       [252:0]  mdsMatrix_32_8;
  wire       [254:0]  mdsMatrix_33_0;
  wire       [252:0]  mdsMatrix_33_1;
  wire       [252:0]  mdsMatrix_33_2;
  wire       [246:0]  mdsMatrix_33_3;
  wire       [254:0]  mdsMatrix_33_4;
  wire       [252:0]  mdsMatrix_33_5;
  wire       [252:0]  mdsMatrix_33_6;
  wire       [254:0]  mdsMatrix_33_7;
  wire       [252:0]  mdsMatrix_33_8;
  wire       [254:0]  mdsMatrix_34_0;
  wire       [254:0]  mdsMatrix_34_1;
  wire       [254:0]  mdsMatrix_34_2;
  wire       [254:0]  mdsMatrix_34_3;
  wire       [254:0]  mdsMatrix_34_4;
  wire       [254:0]  mdsMatrix_34_5;
  wire       [254:0]  mdsMatrix_34_6;
  wire       [254:0]  mdsMatrix_34_7;
  wire       [254:0]  mdsMatrix_34_8;
  wire       [254:0]  mdsMatrix_35_0;
  wire       [253:0]  mdsMatrix_35_1;
  wire       [254:0]  mdsMatrix_35_2;
  wire       [247:0]  mdsMatrix_35_3;
  wire       [254:0]  mdsMatrix_35_4;
  wire       [254:0]  mdsMatrix_35_5;
  wire       [253:0]  mdsMatrix_35_6;
  wire       [254:0]  mdsMatrix_35_7;
  wire       [251:0]  mdsMatrix_35_8;
  wire       [254:0]  mdsMatrix_36_0;
  wire       [254:0]  mdsMatrix_36_1;
  wire       [253:0]  mdsMatrix_36_2;
  wire       [253:0]  mdsMatrix_36_3;
  wire       [252:0]  mdsMatrix_36_4;
  wire       [252:0]  mdsMatrix_36_5;
  wire       [253:0]  mdsMatrix_36_6;
  wire       [254:0]  mdsMatrix_36_7;
  wire       [252:0]  mdsMatrix_36_8;
  wire       [254:0]  mdsMatrix_37_0;
  wire       [252:0]  mdsMatrix_37_1;
  wire       [253:0]  mdsMatrix_37_2;
  wire       [254:0]  mdsMatrix_37_3;
  wire       [253:0]  mdsMatrix_37_4;
  wire       [254:0]  mdsMatrix_37_5;
  wire       [252:0]  mdsMatrix_37_6;
  wire       [254:0]  mdsMatrix_37_7;
  wire       [254:0]  mdsMatrix_37_8;
  wire       [254:0]  mdsMatrix_38_0;
  wire       [246:0]  mdsMatrix_38_1;
  wire       [253:0]  mdsMatrix_38_2;
  wire       [254:0]  mdsMatrix_38_3;
  wire       [253:0]  mdsMatrix_38_4;
  wire       [254:0]  mdsMatrix_38_5;
  wire       [254:0]  mdsMatrix_38_6;
  wire       [254:0]  mdsMatrix_38_7;
  wire       [253:0]  mdsMatrix_38_8;
  wire       [254:0]  mdsMatrix_39_0;
  wire       [254:0]  mdsMatrix_39_1;
  wire       [254:0]  mdsMatrix_39_2;
  wire       [248:0]  mdsMatrix_39_3;
  wire       [253:0]  mdsMatrix_39_4;
  wire       [254:0]  mdsMatrix_39_5;
  wire       [254:0]  mdsMatrix_39_6;
  wire       [254:0]  mdsMatrix_39_7;
  wire       [250:0]  mdsMatrix_39_8;
  wire       [254:0]  mdsMatrix_40_0;
  wire       [253:0]  mdsMatrix_40_1;
  wire       [252:0]  mdsMatrix_40_2;
  wire       [253:0]  mdsMatrix_40_3;
  wire       [252:0]  mdsMatrix_40_4;
  wire       [254:0]  mdsMatrix_40_5;
  wire       [252:0]  mdsMatrix_40_6;
  wire       [254:0]  mdsMatrix_40_7;
  wire       [254:0]  mdsMatrix_40_8;
  wire       [254:0]  mdsMatrix_41_0;
  wire       [249:0]  mdsMatrix_41_1;
  wire       [253:0]  mdsMatrix_41_2;
  wire       [254:0]  mdsMatrix_41_3;
  wire       [253:0]  mdsMatrix_41_4;
  wire       [254:0]  mdsMatrix_41_5;
  wire       [252:0]  mdsMatrix_41_6;
  wire       [252:0]  mdsMatrix_41_7;
  wire       [254:0]  mdsMatrix_41_8;
  wire       [254:0]  mdsMatrix_42_0;
  wire       [253:0]  mdsMatrix_42_1;
  wire       [254:0]  mdsMatrix_42_2;
  wire       [252:0]  mdsMatrix_42_3;
  wire       [253:0]  mdsMatrix_42_4;
  wire       [252:0]  mdsMatrix_42_5;
  wire       [254:0]  mdsMatrix_42_6;
  wire       [254:0]  mdsMatrix_42_7;
  wire       [251:0]  mdsMatrix_42_8;
  wire       [254:0]  mdsMatrix_43_0;
  wire       [254:0]  mdsMatrix_43_1;
  wire       [254:0]  mdsMatrix_43_2;
  wire       [253:0]  mdsMatrix_43_3;
  wire       [254:0]  mdsMatrix_43_4;
  wire       [251:0]  mdsMatrix_43_5;
  wire       [254:0]  mdsMatrix_43_6;
  wire       [251:0]  mdsMatrix_43_7;
  wire       [254:0]  mdsMatrix_43_8;
  wire       [254:0]  mdsMatrix_44_0;
  wire       [253:0]  mdsMatrix_44_1;
  wire       [254:0]  mdsMatrix_44_2;
  wire       [254:0]  mdsMatrix_44_3;
  wire       [253:0]  mdsMatrix_44_4;
  wire       [254:0]  mdsMatrix_44_5;
  wire       [252:0]  mdsMatrix_44_6;
  wire       [254:0]  mdsMatrix_44_7;
  wire       [254:0]  mdsMatrix_44_8;
  wire       [254:0]  mdsMatrix_45_0;
  wire       [254:0]  mdsMatrix_45_1;
  wire       [254:0]  mdsMatrix_45_2;
  wire       [254:0]  mdsMatrix_45_3;
  wire       [249:0]  mdsMatrix_45_4;
  wire       [251:0]  mdsMatrix_45_5;
  wire       [252:0]  mdsMatrix_45_6;
  wire       [251:0]  mdsMatrix_45_7;
  wire       [254:0]  mdsMatrix_45_8;
  wire       [254:0]  mdsMatrix_46_0;
  wire       [250:0]  mdsMatrix_46_1;
  wire       [254:0]  mdsMatrix_46_2;
  wire       [254:0]  mdsMatrix_46_3;
  wire       [254:0]  mdsMatrix_46_4;
  wire       [254:0]  mdsMatrix_46_5;
  wire       [253:0]  mdsMatrix_46_6;
  wire       [254:0]  mdsMatrix_46_7;
  wire       [253:0]  mdsMatrix_46_8;
  wire       [254:0]  mdsMatrix_47_0;
  wire       [253:0]  mdsMatrix_47_1;
  wire       [254:0]  mdsMatrix_47_2;
  wire       [254:0]  mdsMatrix_47_3;
  wire       [252:0]  mdsMatrix_47_4;
  wire       [254:0]  mdsMatrix_47_5;
  wire       [254:0]  mdsMatrix_47_6;
  wire       [253:0]  mdsMatrix_47_7;
  wire       [254:0]  mdsMatrix_47_8;
  wire       [254:0]  mdsMatrix_48_0;
  wire       [254:0]  mdsMatrix_48_1;
  wire       [252:0]  mdsMatrix_48_2;
  wire       [254:0]  mdsMatrix_48_3;
  wire       [253:0]  mdsMatrix_48_4;
  wire       [252:0]  mdsMatrix_48_5;
  wire       [254:0]  mdsMatrix_48_6;
  wire       [254:0]  mdsMatrix_48_7;
  wire       [254:0]  mdsMatrix_48_8;
  wire       [254:0]  mdsMatrix_49_0;
  wire       [249:0]  mdsMatrix_49_1;
  wire       [254:0]  mdsMatrix_49_2;
  wire       [248:0]  mdsMatrix_49_3;
  wire       [253:0]  mdsMatrix_49_4;
  wire       [253:0]  mdsMatrix_49_5;
  wire       [254:0]  mdsMatrix_49_6;
  wire       [254:0]  mdsMatrix_49_7;
  wire       [252:0]  mdsMatrix_49_8;
  wire       [254:0]  mdsMatrix_50_0;
  wire       [252:0]  mdsMatrix_50_1;
  wire       [252:0]  mdsMatrix_50_2;
  wire       [253:0]  mdsMatrix_50_3;
  wire       [250:0]  mdsMatrix_50_4;
  wire       [252:0]  mdsMatrix_50_5;
  wire       [253:0]  mdsMatrix_50_6;
  wire       [254:0]  mdsMatrix_50_7;
  wire       [251:0]  mdsMatrix_50_8;
  wire       [254:0]  mdsMatrix_51_0;
  wire       [252:0]  mdsMatrix_51_1;
  wire       [254:0]  mdsMatrix_51_2;
  wire       [253:0]  mdsMatrix_51_3;
  wire       [253:0]  mdsMatrix_51_4;
  wire       [252:0]  mdsMatrix_51_5;
  wire       [254:0]  mdsMatrix_51_6;
  wire       [254:0]  mdsMatrix_51_7;
  wire       [254:0]  mdsMatrix_51_8;
  wire       [254:0]  mdsMatrix_52_0;
  wire       [254:0]  mdsMatrix_52_1;
  wire       [254:0]  mdsMatrix_52_2;
  wire       [254:0]  mdsMatrix_52_3;
  wire       [253:0]  mdsMatrix_52_4;
  wire       [254:0]  mdsMatrix_52_5;
  wire       [254:0]  mdsMatrix_52_6;
  wire       [254:0]  mdsMatrix_52_7;
  wire       [252:0]  mdsMatrix_52_8;
  wire       [254:0]  mdsMatrix_53_0;
  wire       [253:0]  mdsMatrix_53_1;
  wire       [252:0]  mdsMatrix_53_2;
  wire       [254:0]  mdsMatrix_53_3;
  wire       [253:0]  mdsMatrix_53_4;
  wire       [254:0]  mdsMatrix_53_5;
  wire       [253:0]  mdsMatrix_53_6;
  wire       [253:0]  mdsMatrix_53_7;
  wire       [253:0]  mdsMatrix_53_8;
  wire       [254:0]  mdsMatrix_54_0;
  wire       [252:0]  mdsMatrix_54_1;
  wire       [254:0]  mdsMatrix_54_2;
  wire       [254:0]  mdsMatrix_54_3;
  wire       [254:0]  mdsMatrix_54_4;
  wire       [253:0]  mdsMatrix_54_5;
  wire       [254:0]  mdsMatrix_54_6;
  wire       [252:0]  mdsMatrix_54_7;
  wire       [253:0]  mdsMatrix_54_8;
  wire       [254:0]  mdsMatrix_55_0;
  wire       [251:0]  mdsMatrix_55_1;
  wire       [251:0]  mdsMatrix_55_2;
  wire       [254:0]  mdsMatrix_55_3;
  wire       [254:0]  mdsMatrix_55_4;
  wire       [254:0]  mdsMatrix_55_5;
  wire       [254:0]  mdsMatrix_55_6;
  wire       [254:0]  mdsMatrix_55_7;
  wire       [254:0]  mdsMatrix_55_8;
  wire       [254:0]  mdsMatrix_56_0;
  wire       [249:0]  mdsMatrix_56_1;
  wire       [253:0]  mdsMatrix_56_2;
  wire       [254:0]  mdsMatrix_56_3;
  wire       [254:0]  mdsMatrix_56_4;
  wire       [253:0]  mdsMatrix_56_5;
  wire       [254:0]  mdsMatrix_56_6;
  wire       [252:0]  mdsMatrix_56_7;
  wire       [253:0]  mdsMatrix_56_8;
  wire       [5:0]    tempAddrVec_0;
  wire       [5:0]    tempAddrVec_1;
  wire       [5:0]    tempAddrVec_2;
  wire       [5:0]    tempAddrVec_3;
  wire       [5:0]    tempAddrVec_4;
  wire       [5:0]    tempAddrVec_5;
  wire       [5:0]    tempAddrVec_6;
  wire       [5:0]    tempAddrVec_7;
  wire       [5:0]    tempAddrVec_8;
  reg        [5:0]    io_addr_regNext;
  reg        [5:0]    io_addr_regNext_1;
  reg        [5:0]    io_addr_regNext_2;
  reg        [5:0]    io_addr_regNext_3;
  reg        [5:0]    io_addr_regNext_4;
  reg        [5:0]    io_addr_regNext_5;
  reg        [5:0]    io_addr_regNext_6;
  reg        [5:0]    io_addr_regNext_7;
  reg        [5:0]    io_addr_regNext_8;
  reg [254:0] mdsMem_0 [0:56];
  reg [254:0] mdsMem_1 [0:56];
  reg [254:0] mdsMem_2 [0:56];
  reg [254:0] mdsMem_3 [0:56];
  reg [254:0] mdsMem_4 [0:56];
  reg [254:0] mdsMem_5 [0:56];
  reg [254:0] mdsMem_6 [0:56];
  reg [254:0] mdsMem_7 [0:56];
  reg [254:0] mdsMem_8 [0:56];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  assign _zz_io_data_5 = 1'b1;
  assign _zz_io_data_6 = 1'b1;
  assign _zz_io_data_7 = 1'b1;
  assign _zz_io_data_8 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_24_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_24_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_24_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_24_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_24_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_24_mdsMem_5.bin",mdsMem_5);
  end
  always @(posedge clk) begin
    if(_zz_io_data_5) begin
      _zz_mdsMem_5_port0 <= mdsMem_5[tempAddrVec_5];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_24_mdsMem_6.bin",mdsMem_6);
  end
  always @(posedge clk) begin
    if(_zz_io_data_6) begin
      _zz_mdsMem_6_port0 <= mdsMem_6[tempAddrVec_6];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_24_mdsMem_7.bin",mdsMem_7);
  end
  always @(posedge clk) begin
    if(_zz_io_data_7) begin
      _zz_mdsMem_7_port0 <= mdsMem_7[tempAddrVec_7];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_24_mdsMem_8.bin",mdsMem_8);
  end
  always @(posedge clk) begin
    if(_zz_io_data_8) begin
      _zz_mdsMem_8_port0 <= mdsMem_8[tempAddrVec_8];
    end
  end

  assign mdsMatrix_0_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_0_1 = 252'he2ae70deaf0c8cf495c39e3fea5527947bcbcb4711b0203b1b4c4fc28ced7e3;
  assign mdsMatrix_0_2 = 254'h2071ef6384842615d6e204adaa74831ca1425441a96232b037cfb1cc39c08e9d;
  assign mdsMatrix_0_3 = 253'h16b5fcc072323ce348923b44ff74652f572255c56fc01cef0305f5e6f9a57273;
  assign mdsMatrix_0_4 = 254'h31204f9c18d4b80890a53f812cb40e33ab550c3534b7a9887684919c7389bfea;
  assign mdsMatrix_0_5 = 254'h254c04b40bc3eadd333eccc13ba37693a540e89c55f767d2fb60445c7ec87666;
  assign mdsMatrix_0_6 = 253'h1a62b7b1116f36f33721cd9785817e5abce30102a7da417f602ff3ab4132b6af;
  assign mdsMatrix_0_7 = 255'h5062382a43d09bde7d89f15c20d0bd4d6381191b3ebea8176bc8b7d7d692a7bc;
  assign mdsMatrix_0_8 = 252'h95ddd819505637cb96c616b1ed4ed0f309fa37b03892162dc790c668c477f11;
  assign mdsMatrix_1_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_1_1 = 255'h6f4f19b743056ccde8f99f597612df5e859e5aa7ad726bd061ef82e159dcfd79;
  assign mdsMatrix_1_2 = 255'h6b9ad26fd026137060eea788877cca918bfc02faca0548243449004d083680ae;
  assign mdsMatrix_1_3 = 255'h58d63a324cc98ec7459ebf09a62e67409ce434cffcc1dd7fb3a47213c946e1cb;
  assign mdsMatrix_1_4 = 255'h45f2fae4d13ee525292ae79b9959f91ba286ef3306f5658296f188f707293163;
  assign mdsMatrix_1_5 = 251'h6cb381ba62d1ee1ac93af3b4f917d218ab6a56592fa863063ab78119280584c;
  assign mdsMatrix_1_6 = 255'h5240f0d16b9feb9afde0ae9b805a05a2cd9ec0345182b857bf176846d6092c7a;
  assign mdsMatrix_1_7 = 253'h184124ca691099536c4ab6d3e9f77f9604f8f6b2aab38b770e4273ad19acb0cc;
  assign mdsMatrix_1_8 = 253'h1dc2a509ce49821064065794a0664dd7538e3ea42860b13aadef5c84e0e0841a;
  assign mdsMatrix_2_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_2_1 = 254'h3022b2f2c9ab9fc411561bf52023f21b58956e31550240eb4e9dc4600e4dbdd7;
  assign mdsMatrix_2_2 = 253'h1dc2201448c5103bfb419b288a8387d331c70414a3ca59ae0291d91a31b90570;
  assign mdsMatrix_2_3 = 255'h51042a1ce77e55c544bdad9801ae063654966ce2d257f356ee51d2eed0bbd400;
  assign mdsMatrix_2_4 = 254'h2afc4bfd99265e255120467aef660195cbad68f56aea6f7ea41f5c7ee33363ca;
  assign mdsMatrix_2_5 = 254'h3e837954459dcf257cfdf41c6d005cbc7a61725668af7f82df90396d3c6b48d4;
  assign mdsMatrix_2_6 = 255'h58e523773188da618936eb4f8f1433da7fbd0dbd0f925248139c4f9c053b5a8b;
  assign mdsMatrix_2_7 = 254'h26504905613ab805236818794d0b398c4ddaec7e43711cfb910cf63e7d4f7ecb;
  assign mdsMatrix_2_8 = 255'h4b889b8554199f0382f0658ad5be5c9d0cab0fe7c64f87de667ba03042bcae89;
  assign mdsMatrix_3_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_3_1 = 255'h491fb2665855bb7c2f76e4adfdc5e76e8a1c01eb0a6df858f50ecabea2c0fdc0;
  assign mdsMatrix_3_2 = 254'h3acc493b52d64320c29ad0361fd14538cc0366714c110e7611263573f4a578f8;
  assign mdsMatrix_3_3 = 255'h50dee13f485a92db08746684de5a72fe03f15fdfa99e21919c103a69c6441a33;
  assign mdsMatrix_3_4 = 253'h1536f16109432f8b415dcdff616fc00e37d6f9c8118e091b033181b80db75e09;
  assign mdsMatrix_3_5 = 255'h68ecd80deca2a1f8bc0fdcf71cf0a8174fd9853bbfbf5fd4299429c4adfcb677;
  assign mdsMatrix_3_6 = 254'h2825b745c67751e246041c58916781fb943f272bc85e4437d85b903b38493272;
  assign mdsMatrix_3_7 = 254'h3ed433d6792ba2ab655949fa3325aff66e998fc4fd3d7618b49555c24b82c7e0;
  assign mdsMatrix_3_8 = 255'h73c1f0d1acad8ef465ebc07dc713b280030c8b134db07fbc1e310d1fee1d03ee;
  assign mdsMatrix_4_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_4_1 = 255'h49abe03532aa1c14168039764463f42a85f60ddb871f9f7091c802fbd860b5d6;
  assign mdsMatrix_4_2 = 255'h410b8bdfc4e0a1c1af990ef2c56d018444497b615d67de382430b6333524943f;
  assign mdsMatrix_4_3 = 255'h600c6eed81aba7768b40b10b16d830edd020f13269a15fe515982127abbdccbb;
  assign mdsMatrix_4_4 = 255'h4c15105bf82b305bd1f11972340d5aaea2d0df289e7a0171e3c52bac36216684;
  assign mdsMatrix_4_5 = 253'h17d83375452db559b0171cea90b484868ed18843884be00b72a251e6eaa73612;
  assign mdsMatrix_4_6 = 253'h17cb0bed97766b97efee72aa24e1645b9aa4fc357c23fa624b99ea27d788a1c9;
  assign mdsMatrix_4_7 = 251'h5fc0e35eec4d5046c11c36ea7d0efda3f68a438886bb4f127e47f135110ed6c;
  assign mdsMatrix_4_8 = 255'h592c135482805de35e332277a4cc481e1c0533e770543a3c2a63f64dedab2690;
  assign mdsMatrix_5_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_5_1 = 253'h1ca93da1ac15d8964f26f7b5d3caf9094a402a34d82c446d014ce5323764bb1d;
  assign mdsMatrix_5_2 = 255'h73e5099d4e759abaf77feaae085f7d538835948d3605efc864ae45feb90ed181;
  assign mdsMatrix_5_3 = 255'h4f5f107985e5794b22bb6be4224fe3254f896cff598b6e9062c337f5c49437fb;
  assign mdsMatrix_5_4 = 255'h64755f08d9e027f4e263b939fab3e33fe219448ebc9f1d9368d260512c3731e7;
  assign mdsMatrix_5_5 = 255'h66fe3bdd3b9fffa209fd4764213461888991c94165b879ac08cdbad58b1a5aba;
  assign mdsMatrix_5_6 = 255'h61f7d6875601c29cfe7b19b775b52ba12246f33cb7f5d3b9839572f53a5be7ca;
  assign mdsMatrix_5_7 = 251'h6f002b3ce2d65066d148b29b790496e05f9732fdbed7743d1e71d008c66c75f;
  assign mdsMatrix_5_8 = 255'h4c8122575b4239c7b59c53c46b204e7d5d5b1dad6ef3b9707c9fda7d96dba92d;
  assign mdsMatrix_6_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_6_1 = 254'h3a103844efb5f87d3ab5b262f1ed70a961dcf2eb85204781e20ee0a4bb7bb880;
  assign mdsMatrix_6_2 = 254'h3b122955e7467e0b6b75890efe2865516d1ac099ebb61cf4f4d73699bbafdcae;
  assign mdsMatrix_6_3 = 255'h4ef4b7ccd93c6730dcf6b878d0f8366aed739cb8d38bc6a11f6cbdb116e6ba29;
  assign mdsMatrix_6_4 = 255'h57effae24007bf9a19554415372e60e7595bd64c5f3402d4895d956f05e03e1b;
  assign mdsMatrix_6_5 = 253'h14ef448d358b514bcfbc958565f007d58437f2d5164f712ecb6feab14a8df95c;
  assign mdsMatrix_6_6 = 248'ha9938acc90b69acdbed4cd8d6a48a6ceb6172cf409e931a5405aa7f1fc67e7;
  assign mdsMatrix_6_7 = 255'h5898e12814831b2757c9ffaddf22af6feeba52a6e2bcf1134c28cae78eb709ec;
  assign mdsMatrix_6_8 = 255'h5a09fc4cccbe0bd7bf7d2d6bba7e63ac2c3f7e1c33826939d926001b662a4064;
  assign mdsMatrix_7_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_7_1 = 253'h177ac2d91f98d52aad5752f56498a11db16b3c073d3b19df9fe33064d6fb46a9;
  assign mdsMatrix_7_2 = 255'h649a2eb55182fe35b4921f559d3b936b0fcffbbfd5cae57176070dcb4c25dd64;
  assign mdsMatrix_7_3 = 253'h1f58e70906defe6bfde27f3a0f086229f48e764df84ac245afdfbaeaa76e02af;
  assign mdsMatrix_7_4 = 252'ha40d9f44f38550d7ae7e000f7d1395e1ec6368055b1f73edba0fdb66641b89d;
  assign mdsMatrix_7_5 = 254'h334f359598883584a2c4e0926b6bc6c10773293471288f661253bd15776dc090;
  assign mdsMatrix_7_6 = 254'h2d79ba4b4305359311bded7925d8c8038c6cc2f13500a34acd2e53732fd2c6a0;
  assign mdsMatrix_7_7 = 252'h87be93c95773fafae88fad6122c2be572baea214ac4c78e5aef6df744ed2b5d;
  assign mdsMatrix_7_8 = 253'h1df8bef3816877df6913d93032a3d5d35b79cf0b1c7657d319c0aae9cb57d30c;
  assign mdsMatrix_8_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_8_1 = 255'h67509aa5f56ae1733243a84d0d395f806f2a6866a7d1ce03c1e855d706de42cb;
  assign mdsMatrix_8_2 = 255'h6ea2b5556bcf31b193a902bad23dfa5d592409e88f4b86bc359fab6a31db6bec;
  assign mdsMatrix_8_3 = 254'h3f07f4df1eafa979769e8528a021728ddd99b30e6c8dd6b4760f05dfe54fcfe0;
  assign mdsMatrix_8_4 = 253'h1859cc6783b10c0d759c25c63c28a0e50bc160d4f2728f9c4de5a19a96f7a682;
  assign mdsMatrix_8_5 = 254'h2d20fb3a2f1c0f1f38787b03e5dbee2d16e9571b4170a7d5b96d2835bb950ce3;
  assign mdsMatrix_8_6 = 255'h415fc6edbd998854884eedb07f484aa6aaea42a8c6d72d023404392c4bae473c;
  assign mdsMatrix_8_7 = 253'h16c90e2472ff83f77889f0ff915bcc6c31b182aafd49eabac18f678ecadfaa23;
  assign mdsMatrix_8_8 = 254'h344d280ae7c1c3a31f429ad910fc1df7d8a39e1215e7583549f97abd9b638a67;
  assign mdsMatrix_9_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_9_1 = 252'hba9ecb445146c4959c566070760cc27fe7c097b9460f3baedd80d2a8dfbce8a;
  assign mdsMatrix_9_2 = 254'h32231e920a10b42823b62c2d461da7e4c38d3154d09ff105185a8fd18fd8fd6a;
  assign mdsMatrix_9_3 = 255'h69803a9d27df6188e4901755ea88db87eba260baabfe7f2c466b554c2d137ee2;
  assign mdsMatrix_9_4 = 255'h7213bbcc8b1f96d9dcf92da2243d4b610b092bb0f54114a51e1ee7a4549aeff3;
  assign mdsMatrix_9_5 = 254'h2572fecbc9adba7df2f6b73dc0202ebbe9191b9fdc29dea911726ff2947f80cb;
  assign mdsMatrix_9_6 = 255'h5d55905716612edd129f8bbfca652a51911b1362a41277a294eb62ec3d77a0cc;
  assign mdsMatrix_9_7 = 255'h701d336d3b8b6c99f0364f37a9ac3c279576f3f7a937aa58d0c0ddac05d2a284;
  assign mdsMatrix_9_8 = 254'h2d74ed23d5660c4b04c5174d0ba22944cd0950ecce0fc6a6a2975dcebd54059e;
  assign mdsMatrix_10_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_10_1 = 250'h398dfb3893da73a99d358a55bbd4d3ce5145f9aef57a9b9dff6d3e3b1d5b5b9;
  assign mdsMatrix_10_2 = 255'h4430ffe324fa0cf21864921607d3939320b63017ea897423232e690abb18c388;
  assign mdsMatrix_10_3 = 254'h2717349a1a5b9583266b72767f8c67864ff32de7ddbc009d4d910c23b0c9f9b4;
  assign mdsMatrix_10_4 = 250'h2cd31f77f97844dfc875e590b811fa08cd5068b56c4aabae350dd9df738736e;
  assign mdsMatrix_10_5 = 253'h1c0233c53219c36d2217d1f6022fe0117a873d1a9946e8c79f73451861f9944e;
  assign mdsMatrix_10_6 = 255'h50039822141d582d838e328fb71198b6a7160a0ebde251c3aac1df0755141e30;
  assign mdsMatrix_10_7 = 253'h12fc908af86cc2fb5b9320937b6f2f75ceb9c10e08b55b23320d9c644c50bf5d;
  assign mdsMatrix_10_8 = 253'h19cba5c7b375eb78a1a59de4fac21d9ba560b3d536c5fbadb24749b0fd45fa5a;
  assign mdsMatrix_11_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_11_1 = 252'hf4b668d6fd1a505e46f53f9b633586f8d45710180fabbd3be9fafbee992db58;
  assign mdsMatrix_11_2 = 252'hfbe6b3fe1081abfa0f810dbce2923ccde7bfc66048f78ccf0990d6fbe8415ae;
  assign mdsMatrix_11_3 = 252'hce068ef07eee55c588d18a337b2cf80839d6ccb83bd2a1758a46d973d55a274;
  assign mdsMatrix_11_4 = 255'h705ac9eeffd7887fd3e5ae3e5950570da4c853177d6c52fc4601b1d0bc76c0a2;
  assign mdsMatrix_11_5 = 255'h64f77b0bbacd6d72f7e37d72d2e210d6d3e072110b4dee3d0345fbc0fda3cee2;
  assign mdsMatrix_11_6 = 254'h2dc87c858fc767d189db8b99c2f7d9ac3434641349d0b01d0fd7edcf613cff3e;
  assign mdsMatrix_11_7 = 254'h20668ae74ed8b12ecb2fc6ea77307ed8f886332cea381364a8cb82ca35f56c5f;
  assign mdsMatrix_11_8 = 255'h4f7ea632034a9d837f7291b9790a733063cf77233dfae96f32afdfb24fdf2bd9;
  assign mdsMatrix_12_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_12_1 = 255'h50c17dd204634a8f7a82b11f50c967bb24e68975a185ca8ad8a9e11d45afad2d;
  assign mdsMatrix_12_2 = 253'h1de7b50a9113d25f3d37d0c69faf9eef67901fa05e640e927e4d0caaad4070f8;
  assign mdsMatrix_12_3 = 251'h49c819fa69277315dad164ab598857ba23aa1317d6954b3d945b04f04b1d0d1;
  assign mdsMatrix_12_4 = 253'h13e53e67fc1d184aeb948cc7e076061198288b268c281cfaf0730634b55be7c6;
  assign mdsMatrix_12_5 = 254'h3a7240544240cf9722159162d66b1f7c66c507e13dc0ee8ee8bd7156ff60ab07;
  assign mdsMatrix_12_6 = 255'h4f244140ef8b6a3753be225ae3de29a585d36b7422561c6c8c43dd48c340b9a5;
  assign mdsMatrix_12_7 = 253'h118b0872d0402e4b29c34761fb14dbdd7ad788d265d128fbe4c8b8fa7573925b;
  assign mdsMatrix_12_8 = 255'h70e168ebcb8993e0f7a82dceb27233dbdd02d73754288048df0fb57079b1c439;
  assign mdsMatrix_13_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_13_1 = 253'h15992c3f577b6b0fb3a3560a9e9907e369bc55d01eaead745f22e76e59f31064;
  assign mdsMatrix_13_2 = 255'h70f4727db4ebdd7f4d7c1c5f1ebf6d64f6ecbbdc8b0cf083ea9b77623fa168e7;
  assign mdsMatrix_13_3 = 250'h362d2bfbb46cac87c1467f9919daa3b0e169273393a073de5166dcfe7d52943;
  assign mdsMatrix_13_4 = 255'h5b7ff98ecb0d3874ba7538a37037d53300844f8f399ec577a480d6c71252cce9;
  assign mdsMatrix_13_5 = 255'h535ecf4ed0e9684710faa9cbdbfd1452411540cedcde128092d72e96e6ced64b;
  assign mdsMatrix_13_6 = 254'h23795202d00466e0a20bb2db50e4bd92d0c5a4f66f45f807f7fdc170c64daf1b;
  assign mdsMatrix_13_7 = 252'hfbbeab2e1246f84baa837c000067fb5e20ba51651efccfa3e8db927c0ac7a22;
  assign mdsMatrix_13_8 = 254'h23ac27038c18922b1256276bcccab539b12f7a5ec3840f99651155c93f73c32c;
  assign mdsMatrix_14_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_14_1 = 251'h6ed5d70bf00c2fdb861fa5ccbf997d4a298ba686176ae777e5661323541443b;
  assign mdsMatrix_14_2 = 253'h1e89bdb25c97d01c8bbd541e797e88248de7f1f0caa90c5694991289eef2afb7;
  assign mdsMatrix_14_3 = 255'h558a7f128760cf15fc05775ae4ff4f151a760ce204ef97c73f2adf1203edd66b;
  assign mdsMatrix_14_4 = 254'h3a6c7845d83922d0a8fb652ad6444cbe20718c52f69db91ceb9342948e2046eb;
  assign mdsMatrix_14_5 = 254'h3cc141bb9fd8b17ae3525d8246705e10e20c32f13905ce97b46d54828a4c54ab;
  assign mdsMatrix_14_6 = 251'h4ea9ab7ee38ee8f32c929acacfbb66c6dd5ac3a889cf6c88e8db6235c3881e9;
  assign mdsMatrix_14_7 = 255'h47d766d5111439ef5d50a020c48003ab2e33843a339bf45ce26fda63f08893ec;
  assign mdsMatrix_14_8 = 255'h6a45c745b7cc97d4d5d2a0b84b20653879791564c0c065b096a8da91dc54f0a3;
  assign mdsMatrix_15_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_15_1 = 255'h59eb5ea06d24916a94683cd43b9f7167d4e376ace6428d9b3c1a403c9b561370;
  assign mdsMatrix_15_2 = 252'h9811baeb4619b076bf1ef08d0965a43c306232be4fde95b7a8f46fc65bb8a9e;
  assign mdsMatrix_15_3 = 255'h40e05b03f49f05aee812da4d675bf471f97c4d6cb05f750764c73a63da1157b3;
  assign mdsMatrix_15_4 = 254'h2ae6119b16b1224e144ab840713380c2ae3020cea83fd62254a698e8900bc249;
  assign mdsMatrix_15_5 = 253'h1c0b177c9c714b2f4f46ef9cbb3bf073b79f01d3a9963cf7416a26313a77c2f4;
  assign mdsMatrix_15_6 = 254'h275739c1d93d76bb3c78bedad586e04ff0fdbfad56ef9bc0c4d170427965b443;
  assign mdsMatrix_15_7 = 255'h5e6bfdac5750988e1a66c52bda10eed09ec4703c351b6291c871dc6ab209d1f9;
  assign mdsMatrix_15_8 = 255'h6a160085e96c2a9e3cadbf6160083c19d1d6ce813f83e61202ac9cabf973697c;
  assign mdsMatrix_16_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_16_1 = 255'h516cdaa2ad92dbd4fa34e1287d4a26fffd32d727865b18365839285326212efb;
  assign mdsMatrix_16_2 = 255'h4278a16506fe1670773dca5afd80a75158351142ba2996bb9951212da9863882;
  assign mdsMatrix_16_3 = 255'h5421f6b86837c739c5c526087c43e1eb7063b52ef58250f911cd38b25273a370;
  assign mdsMatrix_16_4 = 254'h2aca81495bfef679abd34df378c0a01ef90b8c93921db699eea172d1e0197d46;
  assign mdsMatrix_16_5 = 254'h200c98ec99262a4ad04fd5521d3df632558e14850bd65ef2dc56ec54f9d9c9e0;
  assign mdsMatrix_16_6 = 255'h6a0997aab038127c86d6c0f2fc9dd3007bd125e369508f1d13135ace136a9d0f;
  assign mdsMatrix_16_7 = 255'h713e9fbfb73ab9a0fe0b313624d88115ebd05c4534b965c079f7ce8d9019349a;
  assign mdsMatrix_16_8 = 254'h3890f1791d91d38eab4230c198b1bab5adf5560ac27193c4b79346ecdc562458;
  assign mdsMatrix_17_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_17_1 = 254'h3af8185151e3adab4385c18ecc00b71f62f20a1a1568ec171c36f1396f8ab171;
  assign mdsMatrix_17_2 = 255'h5975efe15ce1c284166761eab2e9abd9e1b57d772850e82aec073ee818cc0a4d;
  assign mdsMatrix_17_3 = 253'h11fd435cfad0624c339faece569764a4ee7ede8766ecbdbe279208948c553393;
  assign mdsMatrix_17_4 = 254'h350a491b8439c15dcae185482ae9f6b3d9ea9277833ae30066200e6e89466532;
  assign mdsMatrix_17_5 = 254'h2a4da2c18769894e5dd2f46c24ff2157a46b5eea06ae4ab87371851fcb8473de;
  assign mdsMatrix_17_6 = 254'h2f94d4d24ae44df4943ca161198d42f6ff226399699d48c90e9c9e743c0d2f63;
  assign mdsMatrix_17_7 = 252'hc350dbfb61873fb28c45b469cbb2aeb082d23fb11ab708724589c74f5fdf450;
  assign mdsMatrix_17_8 = 253'h1278e0dbc25ff06d2e31cd5d5c07fc22bb1643d90843005026579d4497764b18;
  assign mdsMatrix_18_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_18_1 = 254'h3ef0214597383b1dae1d5a4764f82530654cbf42c06476ab6d91db4137a12fda;
  assign mdsMatrix_18_2 = 251'h636ce1dbf6689aa60ae4d1c50ff505bbe6a985fbf3525585718875f8b1ea84b;
  assign mdsMatrix_18_3 = 255'h52e7b4cc87aa6f9512e22284a92b17d124d5a28d6b247ac8281bff1e46269da2;
  assign mdsMatrix_18_4 = 251'h783284284d4b7e7f9eb13eb79f759a781ff64e484a54367adaacb70ded864de;
  assign mdsMatrix_18_5 = 255'h69634b98d306e0df7269773cabb18fe2c6a1d2ae6f65bd050dbf2862e5cd4e4a;
  assign mdsMatrix_18_6 = 255'h46442d147ef9e77fff91f488b5c040eb47964b52b385f1cd8ac4ecdf609e65a2;
  assign mdsMatrix_18_7 = 252'hf01d1c6f3db0f7da9acf4baa2e0a9f72684aee596cb4cf461540ee785987fae;
  assign mdsMatrix_18_8 = 255'h6a86d4a527b00a9f9c4597559f3fe2b16cdd2d927d92df5bcd17caf428c07c58;
  assign mdsMatrix_19_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_19_1 = 249'h1b1872107c0887ec3bebd020fa27ae4ecb0d89bdf0b057a9c876996d81b7554;
  assign mdsMatrix_19_2 = 252'h87d8578994bf21e0dea1bf9b79a5a2fd7b84eb0eac02b2661dab6e11ff18b5f;
  assign mdsMatrix_19_3 = 252'hb7a14bddaa8be85d7752e01ea04651080b5cf0f133d6c5187845f6eed1cb0af;
  assign mdsMatrix_19_4 = 254'h201ef93b07c416e357783bcd4d27b7a7648c33767a71d30424e20b2368037424;
  assign mdsMatrix_19_5 = 255'h4d5a19f6b87e90d6d1fbb168a5bbe432bf07dbcff620081ac56985853d165ebd;
  assign mdsMatrix_19_6 = 254'h2a4928030e5110a5b93ff892da2e676945a68437d7340eaae4a4dc80856c7d11;
  assign mdsMatrix_19_7 = 255'h6533d6f395c26e6d39441585d7d88ce0d7c7df38300a6e63974595d6fb96d376;
  assign mdsMatrix_19_8 = 254'h299f27dd01762be8a8fc433b3436ed104466aa9167437d5a8d8156ce8fa7ade9;
  assign mdsMatrix_20_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_20_1 = 255'h6779d2c2c5aef13f90093ddcbef36317d72c3d337db1b8f89f1afad2e4ff8c98;
  assign mdsMatrix_20_2 = 255'h5d4ef249e31174be749e340852942e2f1a75289b4665b1397cffcd70a419cb55;
  assign mdsMatrix_20_3 = 254'h280718fb0135626c19c6ecd81f43374fc639217bcdc3485a85e461d0908c668c;
  assign mdsMatrix_20_4 = 255'h4c42e7030232a0733721d85ee94cee73d3b26968f5828db9657010c3bbc35ed0;
  assign mdsMatrix_20_5 = 253'h170f59072c9f4ea4eab2aeeae9047bff333638f80757c8178a5146deb7efa273;
  assign mdsMatrix_20_6 = 255'h631332d64c13fae6e15dac1a918b60da69418fbfcfcf5ee4e463899949e79d93;
  assign mdsMatrix_20_7 = 253'h191dab319fe28d1d33cdb4969faf3ef734d2d86b85a6f0da1eadcc6404e85f46;
  assign mdsMatrix_20_8 = 254'h3deac8c671f0733f1eb7012ce903b3518d815daf9ce584621d8b0c5651064ac9;
  assign mdsMatrix_21_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_21_1 = 255'h5de463161c28fc23f7403743c9adfe72cea7abccc3a3ccded65ef61f9c33d0a7;
  assign mdsMatrix_21_2 = 255'h5698d5cfda1da22a504b1340a083e9fc69b3a1c1187446b3baf513503c2bead7;
  assign mdsMatrix_21_3 = 255'h45d73eb19d17987067f86b47a175f62681ce49d980a6d3afdf5412f033ad8d15;
  assign mdsMatrix_21_4 = 251'h7a5c470422727a69d23ff05bb3a2555949abd601e5ae8b89ed0c9ff15e892c4;
  assign mdsMatrix_21_5 = 253'h18e8029e1f40e7d1ca049135a5540d3faaea5dce7454673efb1e08a0cf5b89f6;
  assign mdsMatrix_21_6 = 254'h380df8f94680cd4dca1dafe448f90843ce87c4b007bd006df6269b4399b835ac;
  assign mdsMatrix_21_7 = 255'h460a996bd67ca01264b0759867d074b67640ab6f3965ab391af881f0611420db;
  assign mdsMatrix_21_8 = 254'h28b1431bc67ab99381339084e6ac1ad14bc206bc33e28b70c6e758c671c3eb61;
  assign mdsMatrix_22_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_22_1 = 252'h97a74133e2ec9a00ee9d54a23a9c3abd2cea3a8440623ed6a5861cbc4e3f431;
  assign mdsMatrix_22_2 = 254'h2e21739eac77c5f55262b38203580735f5f72c590abf0739494739d96f221a81;
  assign mdsMatrix_22_3 = 255'h605a2b136aa3677512c3481129c4aeb52789b08af8c9e51e6e599870ad62a7e2;
  assign mdsMatrix_22_4 = 255'h4e7beec8602762367500465ba07bde6706f2d02b6a2904c2490cc7ffb52b3828;
  assign mdsMatrix_22_5 = 254'h3109dff9cb45bcb264d3c36aa02e17aaee4ddf0918110e2c74273790388baef8;
  assign mdsMatrix_22_6 = 255'h531162294879f0bab5100d4bf588856894f12662568d9b0c360528d55bbe7bc9;
  assign mdsMatrix_22_7 = 252'h808d287b1c991340514afdea4b6590ee8a71acd6d17e80022e55c6f6bff34c0;
  assign mdsMatrix_22_8 = 254'h3f2d4180588ac3bf25ef2b18f522a9b2f551e429325ab3ea6e56cbd77ddf2982;
  assign mdsMatrix_23_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_23_1 = 253'h13f934371635a993e3a578a2e297a8965f4baceb02a2badcb33cbe378b193c0d;
  assign mdsMatrix_23_2 = 253'h17c6a3b48b66d4a91b40172f9ee7f0ada2e90521407e70cb64bf24e32c427324;
  assign mdsMatrix_23_3 = 254'h257221792616867fe5d52c4dee04870dd94ef18a2bd06020e46c68e8cd89aa65;
  assign mdsMatrix_23_4 = 255'h5ce24e1211395223546ae19c3caea0fd946a6c338a512c3b804fa47180d408b1;
  assign mdsMatrix_23_5 = 254'h2df9240a92defc54cb0279fa68333f5ae69f30ec2eefab4a54ff196b4537860f;
  assign mdsMatrix_23_6 = 249'h1ee8dcb2731969bebed19ac7294794a3e09ea6c9bd8cdae60695e204c7f739f;
  assign mdsMatrix_23_7 = 255'h51672d4a8ff7572ba6fd1e79e92428a02932d1fc20da7efbf56afd1d37142f94;
  assign mdsMatrix_23_8 = 255'h6a46d4d08de7866319013ef3524a09cf921a557509dbd4d1de733fb79cb6cd7e;
  assign mdsMatrix_24_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_24_1 = 255'h630b5b287ade824f764734a9ce214a2c3aad6ea3874e53b42ea0712ab5688511;
  assign mdsMatrix_24_2 = 253'h1b8d30ade474e998cc36290a57e97724a92d00235b71666656bda48931a97f90;
  assign mdsMatrix_24_3 = 255'h47520879240ad9753ff670f713ec8a1435c6998ee37ea2de6af27a21edcae52c;
  assign mdsMatrix_24_4 = 253'h13e283ca024ecd99db51102c8e99191dc19826749711d8f4dd94997df1dffa8b;
  assign mdsMatrix_24_5 = 254'h304f955a3b7d0c96787c7e4997be626a1a7199efcb5ef416624206d3e48d3406;
  assign mdsMatrix_24_6 = 255'h464a20f12bc5bfbd79ea4031e245537dbe28ea6bb40b6e83df7e7e83bf2e00e7;
  assign mdsMatrix_24_7 = 251'h610f553854d68fb49cb7ca8c71e5ae1b05c93c15de1f2eef436886b784a9359;
  assign mdsMatrix_24_8 = 255'h60cfecd8f1bd4cd4b7383b41e8f2d1e3e183f0b3e0ceb604b9ed5c0eefe9ec45;
  assign mdsMatrix_25_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_25_1 = 254'h2c640e2ad708601adc094398b29010e97b46bdc8d0aef85eea20a8bc8cf46760;
  assign mdsMatrix_25_2 = 255'h4ed9bee35999d8b2f845ccda02a12d8b8aaa74d53b02f1eafa69105c482ddc7d;
  assign mdsMatrix_25_3 = 254'h21edc8e33853ed4860ab89ed5061e1978a216b5015447115c72d0cea8800df4c;
  assign mdsMatrix_25_4 = 251'h7484e3de35f3a6a15e3d5db788b6b90f428f3f0a155aca173e39d5b67a6069d;
  assign mdsMatrix_25_5 = 255'h4f55e813b57b630ec331bf1dc11ebd262349b2b960af4ee324777f25648bb47a;
  assign mdsMatrix_25_6 = 255'h439baf0316112b8537e4b738889d75ec8eb4d4682862329810849937b9b56037;
  assign mdsMatrix_25_7 = 249'h1e8f9ba8ee65c086fd941709fbbc9b0f9d25857f5ec86f43fb7693d5541ba13;
  assign mdsMatrix_25_8 = 251'h4a3d90712aadbad1eabb88a899efba6659288a60cf3adddabcfd17201ff37cd;
  assign mdsMatrix_26_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_26_1 = 255'h5daab91c7185905c992df95e47882d96366dd51dac9df1cc3ae6574b6a0910b5;
  assign mdsMatrix_26_2 = 255'h5bf07ba9054f7243e9332c356fbde21ec61168336ae73668efbb4ff85822040e;
  assign mdsMatrix_26_3 = 254'h2d7aa479261667a64b842bcd53c377b122017a2ec6cf5028ee3f413a656ca9ac;
  assign mdsMatrix_26_4 = 255'h50d6d89bb55087b095d5efd9b8452769e088cfe4d4fede0aef04b3c22ab3d19c;
  assign mdsMatrix_26_5 = 255'h63828089c137f35dab8af26aebb5bafe5ab3ca9afd752c1df112bf7a89be37df;
  assign mdsMatrix_26_6 = 250'h23e40b30e972108034240d29e22ac5d7b2d3d21954a8bccc0153e74390364c4;
  assign mdsMatrix_26_7 = 255'h576a96a5df6951c3ddc2eb98ab23f6522a7a3ccf515b99e3e9268edd5771c774;
  assign mdsMatrix_26_8 = 254'h350ca06b96a353fb8282b44809e36c06a4d8394f025cd47b3ea2e63a3c254f8b;
  assign mdsMatrix_27_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_27_1 = 255'h67b13892abf80e7ec7ffd6e92a550a7816c089b39cb8979c17289781b85adb80;
  assign mdsMatrix_27_2 = 253'h12abcb56fd0298cf1bbf62220ba22d84f228cbdc59efeb0ff58544abcb749543;
  assign mdsMatrix_27_3 = 254'h2f0ac4673b6008dfa8d46d9c883d98582ac6d256c56a759225d6bdaa6b668f68;
  assign mdsMatrix_27_4 = 255'h53dd17320bf9b9e2776ba617ea23e85ecbf4cb02957ae0dffe2826c8dc8ce755;
  assign mdsMatrix_27_5 = 253'h1584c09d9321b21c6a8113775ca7150afbea329bd9bc8300c6eb79f63af9759b;
  assign mdsMatrix_27_6 = 248'hed483b89d8a7c74b9cc48a62b8b91e3a25fd149a4ba7c170ead5c66084d201;
  assign mdsMatrix_27_7 = 255'h55c8da3c35a750469eee83001147a4d395d03e819cf3b374c1b272f8892db1e0;
  assign mdsMatrix_27_8 = 254'h25c51ae13be126247bda9db265a57e6d1927055ce4b0d05438a0e03c3c138be4;
  assign mdsMatrix_28_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_28_1 = 255'h5a1580d12207cf9f2be5681cfe55c7549e5fed4a539251f84cf536175fa6abaf;
  assign mdsMatrix_28_2 = 252'h89e436563922d8ed1c90bed26b3b71a1b96aaada1678007e9dbde362efb7dc7;
  assign mdsMatrix_28_3 = 255'h6267edc2a716cde7b11ca2f9cbe5079f412ed865e07bd9024ce894141105ac02;
  assign mdsMatrix_28_4 = 251'h6c7d6fe783efa9f730540b2b7d2b17933c215334633977c21ff9a3728737192;
  assign mdsMatrix_28_5 = 253'h1fbc9e57eca8769acfb22a7921dafbc83ad601ddac022538e92de314c95830e1;
  assign mdsMatrix_28_6 = 255'h54e08437681700e0fdf23f993a4020766cbdcb8eb02099e6b36cbb2d57b210e0;
  assign mdsMatrix_28_7 = 255'h432c0f0c54398ee54438eb5e4c029a326e3f55d37fff0f77e3ccc56d93947993;
  assign mdsMatrix_28_8 = 255'h598e40ba0c3b2a00d83ddcc5b395a6a7ef90432d03fea89a6538a6dffc0e7588;
  assign mdsMatrix_29_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_29_1 = 255'h493e4845ac9f18a95c3bbd29edb40fa2035202c1b45eba690b379fd4b4daa3f2;
  assign mdsMatrix_29_2 = 254'h3219b8efbf2aeade3d0d4cb25a3005aab4ab722f97abc21b78c8f14283947dff;
  assign mdsMatrix_29_3 = 250'h3c30c7ab0a0618bc590d297e7321fb6964f3b611a9c2c59aa7f0f38e2b44257;
  assign mdsMatrix_29_4 = 255'h42f687a064a1aeaf9d5256a4e97b860877376cfd376cfe389724ed92590feba5;
  assign mdsMatrix_29_5 = 255'h5bd649b4c7477bb3524aa8d89e91cf4c994c8c06711b448c91025ad102f702db;
  assign mdsMatrix_29_6 = 255'h66d4a7e2b0e89a928b1cfd11640237bfd0db3f5668a42eb9eae8fdb5c54b4523;
  assign mdsMatrix_29_7 = 255'h5ad1f6743f82372a0862f95ce6ec1459d138be5f21a81c8542093817fdef0343;
  assign mdsMatrix_29_8 = 254'h37523c221ddb12656bb29710d8706b923400a82324f156264bdf8361206d63a3;
  assign mdsMatrix_30_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_30_1 = 252'h9e7d0115a7c77a75c331cb447e4c089ceba669765b8307862190a7a1c24f033;
  assign mdsMatrix_30_2 = 251'h598e4b4b7fdb301c6ccc4f131fd804d62af67c7d0e40d5d9572d36c5f035563;
  assign mdsMatrix_30_3 = 253'h10ba2f4adf6c12033f33fbdeb1e03034cfdad061fca20d1c7e068755496ee47f;
  assign mdsMatrix_30_4 = 255'h5402c777600369a94c62ebe78eda6495405e4964725a2265f22fcaf7a454f732;
  assign mdsMatrix_30_5 = 253'h1be7d227baf859535fedb816a807082b4116fe3f8ad46fd6c529b4d68bae8498;
  assign mdsMatrix_30_6 = 255'h6bec27bf95650a2145204dc0999b369b008465ba6f77e5a4a6531ef667025d6a;
  assign mdsMatrix_30_7 = 255'h64b99677990cc9eaacea8e39e922e16bad3e50b26f6c63dbb2c2e6716b30ce9e;
  assign mdsMatrix_30_8 = 252'hf4b374aabae772f73e55361384bb3379b5dc99f220954b9b90221bbd97ba3a9;
  assign mdsMatrix_31_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_31_1 = 255'h59330f88e198af3c54ba2623585313084893404302975098b47821b607a83339;
  assign mdsMatrix_31_2 = 255'h42b66a24336b01725a55dded9f28a9ed65006cd398bc27aa16ea34e87ad00874;
  assign mdsMatrix_31_3 = 252'hb9a17c491f56aa9763d377cf59d5a034c23548e2bb914ac71deba25f682590f;
  assign mdsMatrix_31_4 = 255'h401e3cfb427614d59ff1cb8677da28645884d75abd02b7e3e4b1f2c8263b3287;
  assign mdsMatrix_31_5 = 254'h312ba5b476e51066b61e0b15902f7a1f97cce785b3d3f89a5cca5f9486dcf363;
  assign mdsMatrix_31_6 = 255'h64258d9b7cfbf55a7f051042c65c2b638be925dc839f32a4c1d8beabbef27918;
  assign mdsMatrix_31_7 = 254'h363bd29b8d18cf12706aee676f71790303c590545bb63c5e42a5e79e02cb6bce;
  assign mdsMatrix_31_8 = 254'h285550d9e82d3eb338f4426bf918e263a8bb0ad340ffc5e6c7484db80c268c65;
  assign mdsMatrix_32_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_32_1 = 255'h41b77b0358b8c007004df3c7f0eb57fd3bcbc59e057f27c16092be13bdd34847;
  assign mdsMatrix_32_2 = 255'h6f3eee4b6e66c2ac2d4476c142a3128bc992689d92aa4a5efa4287ed78028e3f;
  assign mdsMatrix_32_3 = 255'h534d4535a18e0f6abd559c4b8d642b2245e8c2441fccde3010c8dea7715cd912;
  assign mdsMatrix_32_4 = 249'h12144ff0e6f092b79473d6225cdebbff805aa3c59c017e142d60978c8687eef;
  assign mdsMatrix_32_5 = 252'h8d2c9b898f6555091a2b3c270ce2a4a6f8c44c16e195d471631c5931632245d;
  assign mdsMatrix_32_6 = 255'h4d2ff81e7aa39fc18989b261ab87a17104c245aef5e26a605027402f7bf9dbe4;
  assign mdsMatrix_32_7 = 254'h2e09a82d3f08299a11ce722e81892911c235497f915e519ce85f8151fc837d40;
  assign mdsMatrix_32_8 = 253'h1b2fd4c28cb4def06587bc7e9c50c120525ed166a8c286614622a8b0ab46b508;
  assign mdsMatrix_33_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_33_1 = 253'h1fb8f41fac3e9ada0bee572c3c582dd8b0da2b5cff12cbefb5e3a53e1e6d875f;
  assign mdsMatrix_33_2 = 253'h10fa891630ca78b7286fd1c1170318494777f9e03e8a74ed2306514510cb7724;
  assign mdsMatrix_33_3 = 247'h779bcdaa766cf8c0db497fff07a3176d6bf6a3342178022d9d7b09b4d6323e;
  assign mdsMatrix_33_4 = 255'h5d3f065d4758140b178f0e413dcdbc9057a8828dcabb60387584d7991b121c32;
  assign mdsMatrix_33_5 = 253'h16f0673125005db778a13c5937e44fc0af5274597e5fdfefc0c0a61a609be8ec;
  assign mdsMatrix_33_6 = 253'h1045428864505829e7b8983b75ecffd333db7d77c275684488efb5791a508ccb;
  assign mdsMatrix_33_7 = 255'h6f3cef1bf02ea87c495b724dbc24465d0bca98b27f940af5ac092075aeec1567;
  assign mdsMatrix_33_8 = 253'h104317ba1487f1162f6282a1f2fb118e2689ab2a5c516c20d2392cce398d98fa;
  assign mdsMatrix_34_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_34_1 = 255'h66516e291b6904ec8a91ff62d3d3679da43cfcf063d8c6dab3bea876ffd6ad26;
  assign mdsMatrix_34_2 = 255'h69942af62734dcca96393c9040a7059e0e046810a66969e63307532e2e99662d;
  assign mdsMatrix_34_3 = 255'h46572881b8d794716fddd089ca9012d19e04aad8e93727445c15e0058abd6474;
  assign mdsMatrix_34_4 = 255'h637ca81c1dbc15cb3ff1503b7c1aae01f989937a9336aedf0d5dd93ea85ba695;
  assign mdsMatrix_34_5 = 255'h4321b11c6384dacc0fd898b0e94449ac52e0009da8e1723300dcc62ba7d415ae;
  assign mdsMatrix_34_6 = 255'h519fa79dccaa43e69d73dbd52064cc3faf34d09cec637c9b84f86c8f105b4585;
  assign mdsMatrix_34_7 = 255'h5c42dd52953efaaee5ce39cc5e274119ab05746f2126a14363ee85150a38a2e9;
  assign mdsMatrix_34_8 = 255'h5a9599aba98981d74d1bffdfe76b4a49db708d8300ca1f359953ca5518a763b1;
  assign mdsMatrix_35_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_35_1 = 254'h3d6d1ad8691f9dd65b1a79725f6cc4ffd6d9e03c66d5fd1eed9b46e03733c1c7;
  assign mdsMatrix_35_2 = 255'h4fdd586477b705f90f043d3cd719b250acafbe38012a7e71e198f16cafc33a3d;
  assign mdsMatrix_35_3 = 248'h92f76575d223e82d86db4f6d2a47da84d6cadd7de6f7910a95b5d7307ea084;
  assign mdsMatrix_35_4 = 255'h40fc36ba8990575e866b9885f9ea643647c354cd8803a6ecdb663e308bc37dd9;
  assign mdsMatrix_35_5 = 255'h5659e89b5cbfa3e9836ee53c66b055b678b15d8f360f18d236eb8d3bf45a3a69;
  assign mdsMatrix_35_6 = 254'h2c5d4561025c9c2c506e86e810ed8254a8d7452a5cad401c1b48bc5222308a0e;
  assign mdsMatrix_35_7 = 255'h5df3ef1fa1a42c0e59351a29256bcd6fc3150cad3407373ace5417985e4dc98a;
  assign mdsMatrix_35_8 = 252'h8fa225c2d5540f16d7b1aecb73a472879e1eb1b86a6d7d8a5d5b3eea7c25d92;
  assign mdsMatrix_36_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_36_1 = 255'h57fd7aa1c1503b01794c2b358988b8acb35be9fa102c766631fe46287d4d4743;
  assign mdsMatrix_36_2 = 254'h29a4b0075e9611ca4cbcf917a4ccbdf4276e6974062a2a3d50559bf829624242;
  assign mdsMatrix_36_3 = 254'h3fc8119f94c4874af1cdddf6f6e9a6f7b46719aff734bb5c71eb55100ad5a894;
  assign mdsMatrix_36_4 = 253'h163d1c44791f303bae81edeb75fbfdc0a0d492547bc5b6dd9d52cf1e7486aa58;
  assign mdsMatrix_36_5 = 253'h1c7da5d427374811c513fe8b1b02bc940b6cbe41ab0fb070e26008c139c30dd1;
  assign mdsMatrix_36_6 = 254'h3cc803ac0d0d0d117112ccbcb7ba332048807c5c5da1fd8962bef871d115fac9;
  assign mdsMatrix_36_7 = 255'h68727d6fc819816f8a90b4d532c844f921b6619ecaa354f1c6dc8917497e259c;
  assign mdsMatrix_36_8 = 253'h13c4cb6e8409cd3bccc241fd532f3b2d035cfd0459ac31fbc606d6214eee27ac;
  assign mdsMatrix_37_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_37_1 = 253'h1630ecf479ce169fce52d6242d454274fa2c4dee5268a1f42c936cf779743c95;
  assign mdsMatrix_37_2 = 254'h24d7374110e9e8dc9c845819a196551eb537d03472e2c9e6cf3f000690c36a1a;
  assign mdsMatrix_37_3 = 255'h68f30df5827e3cbc579f85deed7507e721c8d41fdf0154ec635c278b0469176f;
  assign mdsMatrix_37_4 = 254'h32d6a8b55b0c3d27195912381978aacb03ee6889f04a44339b2100e3de812cc4;
  assign mdsMatrix_37_5 = 255'h5d0c12d7d8bbeb2e4f6aa44827f261f59e67745c921ae1fee698841e1cd1d175;
  assign mdsMatrix_37_6 = 253'h19933e5df3335cada9a3e1d3515661fcb1bc747fbea150e1dda505c45cc4ba8b;
  assign mdsMatrix_37_7 = 255'h53c970c9652d3399beaccaf700d710740607537b12f32b7565fe50d79c7dcad0;
  assign mdsMatrix_37_8 = 255'h435f09ee3e0c5b45811c1e0106dd51e0354f603b1eee3c5e8ce6a11f50b80b1e;
  assign mdsMatrix_38_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_38_1 = 247'h7075cd3dcabe2681ee0ee1a03dca1dde84ec331c44454ace2e16b369b8008d;
  assign mdsMatrix_38_2 = 254'h202224643e3eb1eeaef43d7d7e68a264bde64a833dc80ece6cd42124a6699c40;
  assign mdsMatrix_38_3 = 255'h5e45f8dc78ec120978c73ee6ce3dd3845eb5634d3606baf02d56cf451f404c81;
  assign mdsMatrix_38_4 = 254'h25d70f3670cd45ffa4e2fe3a2728346bb22856ff17c258fd59c6c682443d62a8;
  assign mdsMatrix_38_5 = 255'h48043039b003a24aa72d91fb327c4801415d41fc145ccf95836a20e46c366711;
  assign mdsMatrix_38_6 = 255'h42f07b39f09a2ca12bc61d22760dd459546cb0fe50ecc591d9bb99cec4b9a046;
  assign mdsMatrix_38_7 = 255'h5235622022fd7eae32eacaaff2dd7a9cb80147f1a5c4bd7369da941fa9d54c44;
  assign mdsMatrix_38_8 = 254'h35942df48aa0fac5d2d697555da04ce51209336a8af6886df183571367442674;
  assign mdsMatrix_39_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_39_1 = 255'h65c49096ac92bb87357b5cd5b23ac5f5bceeb9829ce07740047f733d834eaabc;
  assign mdsMatrix_39_2 = 255'h5f15a1e793f432350f9eeefd325fac7c702aae19e99e60b26ffd06db5b3d141c;
  assign mdsMatrix_39_3 = 249'h13e1a1fe18ac90aff93741ad5fdb640fd26968f7596f8697aa9c5bd7005032b;
  assign mdsMatrix_39_4 = 254'h266d6c295e1a36e9faaea472e1960cf24f2e1ca3b4dee11ba8595935d5704401;
  assign mdsMatrix_39_5 = 255'h59ed3ab71a36589c93456276047aaa6557a02673468ca743ea3529ac6da878ee;
  assign mdsMatrix_39_6 = 255'h641b043257831492670588e8c6411b22e346736af99308dfc992f79fa0698d67;
  assign mdsMatrix_39_7 = 255'h508ebcfbd59eedcd3e953ecc965ff62812536e45644416a898465c7097807e8b;
  assign mdsMatrix_39_8 = 251'h78230dbed2a0742bb0b96185f758ec1b920f00a76d300a6dddb2f65f3fad6b8;
  assign mdsMatrix_40_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_40_1 = 254'h2a4332a43b5be698778ae9e7ba0fcd010d1a4b5d28e4fad748df00407717dffd;
  assign mdsMatrix_40_2 = 253'h13882eb91b6f8e3c93fd919cf9cb893b4a5f794165aad0b31fde6218b0e7d0eb;
  assign mdsMatrix_40_3 = 254'h3872b6efe3259e9e0f3d822be00427d511fc38807c8d0895bb4b91206f05dfd4;
  assign mdsMatrix_40_4 = 253'h149d6026b4ce6af8a3b7afafe6dd4f13987827aaf931aa1bf45bfdfc18947c2b;
  assign mdsMatrix_40_5 = 255'h47c4c086baba1a04b70b6e233081cc72e361616f040f2175c873ab229ff3cd8f;
  assign mdsMatrix_40_6 = 253'h105448e76abb683d0f9cbbcba819a6d18abc8ccc1b3eedfd354c8b08d3d540ec;
  assign mdsMatrix_40_7 = 255'h60cc1fd364c8beeb1b1edfb923919bc389618ba9c6d558102f59d05b2a317c68;
  assign mdsMatrix_40_8 = 255'h50ec4a1234d0114ad980b4e7380194de98046d8049b686ab9e4e3ce55e2c29e3;
  assign mdsMatrix_41_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_41_1 = 250'h203d03330ff01a1412f0ff74bc7ca591e6139c8f2c8f00fe0c274e8ed80107e;
  assign mdsMatrix_41_2 = 254'h2c95ce4bf8b76f3d74af45ced953768c349cb3247f08df045c7b2d214eb035a6;
  assign mdsMatrix_41_3 = 255'h656afc7a265450f5dbf0454c0393e2dbb64327384f5a56e3d7215790c17d35e0;
  assign mdsMatrix_41_4 = 254'h28b56060d5ddb92079bbc79706f84ec3ef2e24ff906c70938dcbf06786f782b7;
  assign mdsMatrix_41_5 = 255'h546f7adbc51b7be1915d5b38d33839e7ca56795395879acbcb06fa6f70a94a67;
  assign mdsMatrix_41_6 = 253'h1dab908f1902b60ca627a6d48807093bc9e19dc4609431ccf34bae9b8f796b75;
  assign mdsMatrix_41_7 = 253'h14f70f2d2101280d22296242062e143aaeecbf910e5d032ef9e8e2c641c03da5;
  assign mdsMatrix_41_8 = 255'h66b2fcce551d7dfc3ba21ffa2b6298a9d287199f8220f0d2e685f20f8b7f2f03;
  assign mdsMatrix_42_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_42_1 = 254'h25aed9ef048f71dd3a9203d19aa2468eb40a3de043065221d2a1effb8ded6dc1;
  assign mdsMatrix_42_2 = 255'h66a2eb56490903d1c7b2b7a0bec3d28152d98a8d6eeedc988b70a633b7118ba8;
  assign mdsMatrix_42_3 = 253'h1b728ec5aecdea64f49b9be969d3b169562dc21e8764e375be349258e5b95611;
  assign mdsMatrix_42_4 = 254'h2aaf91c4f619713c000fb8d0655d2184477939a6c984f692aee7ad23c5dc9789;
  assign mdsMatrix_42_5 = 253'h172768f361a4818cad3c50daee873bd1a410d835096fc79e198cdb86b1fea0ab;
  assign mdsMatrix_42_6 = 255'h6747b6167c6b7a4e6ebbed02dced0ffdc59fc95e3869bd4b9909391045ab0f7e;
  assign mdsMatrix_42_7 = 255'h5532a916738271fd93986e4ef9891c026d368e5ddf865bacacbbaa80b0d79d3a;
  assign mdsMatrix_42_8 = 252'hd36769d57a4b99cac5ce1d7250898e845321ea96889c83d9f3b03ca442d172e;
  assign mdsMatrix_43_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_43_1 = 255'h4a8ae43b670b540dd6c2092283bb6534bbf8c7f8bcecb20c42909fcf12ef6b54;
  assign mdsMatrix_43_2 = 255'h71a27c0c1e92100c459a4d4a4b38c18ddeac3e360fb1ebdf5c1fabaa230e7270;
  assign mdsMatrix_43_3 = 254'h27fb3f08ebe5256fafdccf19d98fa7cd38ae7561c7da0add990fd770685d0a05;
  assign mdsMatrix_43_4 = 255'h424ea6a2d42b91eadc9e7eb2706a1df8cb389082a733bdd458d1c846a53faa01;
  assign mdsMatrix_43_5 = 252'he3f004dd3346aba664f40842f680831ae585787c356fb48ef53422aef108056;
  assign mdsMatrix_43_6 = 255'h4bfeed35e6d6d4e19c23c7f82d0d168b7cb5fb98efda778cc217e4ce62f9a403;
  assign mdsMatrix_43_7 = 252'he98c6d55ffe2bd6959d5df4f4671db6c859b1ccbd6cbe02a078c073e1f70d2d;
  assign mdsMatrix_43_8 = 255'h4d06d586f7192cae889852da1bcdf79e08f6f7f6145040486c026ff82e4b77c0;
  assign mdsMatrix_44_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_44_1 = 254'h3de87296f1f3bace38dabcb0a485afd498fd1e03dd1d7a32512b277c51ca04db;
  assign mdsMatrix_44_2 = 255'h59f4ad12176619df953d846a8924006e1483c202eb383d2108716b20d86dc855;
  assign mdsMatrix_44_3 = 255'h5e7985a43d06556a995e0238f9cc1febef4bcc9e7601a61e64be904a3ebaf0d6;
  assign mdsMatrix_44_4 = 254'h3649a112e088f9cbbe3025a0d7b8b4707284816993368273b1074c7c74a6a670;
  assign mdsMatrix_44_5 = 255'h5276f98e26dc08264b5d781b68db25d3177142a55287e2ea959a2e829b1d5998;
  assign mdsMatrix_44_6 = 253'h1fbc2cd7f27c095f156d015542bf76f8cb732da182913535c190263db7d36836;
  assign mdsMatrix_44_7 = 255'h5dc33a2c010dd2aa98eb17592e136fb9ef40d440f8a131dcba6543d1f1cb4f9f;
  assign mdsMatrix_44_8 = 255'h629ffcff7682e190600707471c73ee9567d5282eeaf7586e8044bd3bb1636b07;
  assign mdsMatrix_45_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_45_1 = 255'h5b420982dfd283f033c33b77a6095b9ed3dba475116d90f3c2e7b54b8651857e;
  assign mdsMatrix_45_2 = 255'h40e0e470bff8b97f52e4ddfe46b0abeb9dbe90dd0e21d6fcf2ff3ea48bddbf1a;
  assign mdsMatrix_45_3 = 255'h6921a6c9273994552564df639521a31af9e020d3e8d919d7ec927b72ff8d47a5;
  assign mdsMatrix_45_4 = 250'h21468e36880ab2a53d511085f9ef0a371fcab207e2ef170cb065e7f305cf51e;
  assign mdsMatrix_45_5 = 252'hfe82f8518027cf7ebee62acecec4dfae44416da0d1f1eb8259c1d696d77d46f;
  assign mdsMatrix_45_6 = 253'h162509b92eb857f3d379d392925c589f02baa2a658be68fabb7441c1de2101fb;
  assign mdsMatrix_45_7 = 252'hbe6596cbe46d363265f0ba65e930e2ee0bffe655a5d0e562daad9eb52520064;
  assign mdsMatrix_45_8 = 255'h47fd7b61c7526f7541d0fda0fc7783c96e3a54c722b307029b95d77e5df48ff3;
  assign mdsMatrix_46_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_46_1 = 251'h4c81f17484ae9af6197461fc0d02d73d763624fecd621f7d91155f492e8a885;
  assign mdsMatrix_46_2 = 255'h602d548a15bb33856499d67327da2a625882aa27e9bf429c070a70f14b95978a;
  assign mdsMatrix_46_3 = 255'h4f4cff3889b4d505d5155e8b1f4eafc6f24e1adba7882c2f0323f53af42c9308;
  assign mdsMatrix_46_4 = 255'h48d36e9e54be7b3557eb3d277b4fca125351e30e390b3ab78de8a523a4606278;
  assign mdsMatrix_46_5 = 255'h5d790b9cb4bf7247499b17a844e2f96e503c21aab7492d941b7303ca4dfbf0b9;
  assign mdsMatrix_46_6 = 254'h3c83a50ae2b33bfb9db4994730845eff74214622eddcd89df2d9b31303513334;
  assign mdsMatrix_46_7 = 255'h5e2d05fd688ce0572c243e91d2562cdcce3161844045cfa06ee11c9b6259f616;
  assign mdsMatrix_46_8 = 254'h35f434fc484fa5941f1a3d4fbd9fc01677a8cae2b16c4aad94bf00d95de37402;
  assign mdsMatrix_47_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_47_1 = 254'h21906fcc59a7e52e42ebf6e1d17802baa1fc0b9bc38fe2f34753aa8aa69a501d;
  assign mdsMatrix_47_2 = 255'h64c5cd31eb2bc73a4aa9a04f65b54b5b74c0c8ea199922e5d77c0a76c8a56354;
  assign mdsMatrix_47_3 = 255'h578563fedf27e93b78298c3d4fd95086cffef5ae60d2b992ab882e3987f0678b;
  assign mdsMatrix_47_4 = 253'h1574eaa64229f844191f83f7d743ce0884756f8cdf2ebc0da887268875f125ab;
  assign mdsMatrix_47_5 = 255'h42884f2645c3f8d51d30acb89900a848cf658bd50d241c834d32f0760a7bc263;
  assign mdsMatrix_47_6 = 255'h645a96745779449cb2c1965a013f03516d0e1d8d3ea02d1cafb417ae1430896f;
  assign mdsMatrix_47_7 = 254'h240332a78cfb5111f01aed34b047b21ddf9bb7060bf503100319499a42a864b7;
  assign mdsMatrix_47_8 = 255'h705a2d7221d521feae9803298a9e5a0abe56f624056e88aac2ecf6fb02a4d7b5;
  assign mdsMatrix_48_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_48_1 = 255'h4cae4938afebdda388dcfc88e9256f35ab7786e3b7501972292749401c87bd8e;
  assign mdsMatrix_48_2 = 253'h1843081dc1ca3dae4d062e6b52a21d5c25178189e6d3131e3c5b819268dc56ff;
  assign mdsMatrix_48_3 = 255'h68ce6f2144d8412885782bc4b5b2cde615f18c6b26928ac6b083aef856c3c739;
  assign mdsMatrix_48_4 = 254'h3c1849efc36e4e5313388f7e886c5928f8013ee1033502a6abaddf11f6fe3612;
  assign mdsMatrix_48_5 = 253'h181675c978c40f5ef3ccdf65b24b6864ff97b9683e9e17d3022c96059ced0761;
  assign mdsMatrix_48_6 = 255'h6507b0267326b24b76ed7cc1f9561cf055e2fc4f331bf50a5e9b69d78cf10b2f;
  assign mdsMatrix_48_7 = 255'h605dc16022a3879d87388b3d8232ce29fcc2114044fcdb259ec161e92d8fb659;
  assign mdsMatrix_48_8 = 255'h70d536ce3bf29f642919bc05c2b6652e7795f58c8e7031f127772a9a61b15bce;
  assign mdsMatrix_49_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_49_1 = 250'h2e2e504bf202a319e1e5c1f9c9a1c54e0b80f7819740909478a6bdb5d0360ff;
  assign mdsMatrix_49_2 = 255'h714bade21b8a79f4b867ff57973621f0c9ccb570ab40624af15aacb22e63fbf4;
  assign mdsMatrix_49_3 = 249'h1f764e34d086cbe14316222aa02da8cbb66957eea23e4992f2b4cb3f7dc047d;
  assign mdsMatrix_49_4 = 254'h22b59b4737e788c6d21f3a4044f990318ac86ca2217d18f2ccd7d555e0f27854;
  assign mdsMatrix_49_5 = 254'h2456e7f11274247d35a48f0dd461819dfe5eacd130a1cf27cfeedbbdd6b41752;
  assign mdsMatrix_49_6 = 255'h708106b193cf43ab305a7855179762d34f8f4f99a26729e7a8d9e44e688e276c;
  assign mdsMatrix_49_7 = 255'h46b2161b1a36332492cdd50b9b4c22ca258ef002845b5a6c8ef359e37972a5cb;
  assign mdsMatrix_49_8 = 253'h1081e33db8feb76617eff224cea841621d048e30f2fa69cdcd2f55ce99195676;
  assign mdsMatrix_50_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_50_1 = 253'h1da6fdad55f423a213e7a6b7bbbb152234294e29474d73475047906dc3a4d425;
  assign mdsMatrix_50_2 = 253'h1331f2800a40b2a9566c87f1aa8ad1f6fe2e30653d8f48026052f8d04ef8e06e;
  assign mdsMatrix_50_3 = 254'h3f21eeb1c255e69ff579835de9ef36c446f8d9996e65e4e27b213a389be3308a;
  assign mdsMatrix_50_4 = 251'h588b1a7422a72c6992ba5caa2158ca5e1c4d9d76bff6e552ab3e6a2dadb8412;
  assign mdsMatrix_50_5 = 253'h1a14984fa528d9a9a532a892c40aa5b04c31527a51143675636b20a810a9e2be;
  assign mdsMatrix_50_6 = 254'h2c49864c6019f93499bc5663e843232562ca80b99202609043e255582ca2db24;
  assign mdsMatrix_50_7 = 255'h479526240b00c65d88c3f0d3939c2bfbdc1552cc9a40555ea2602472607280c1;
  assign mdsMatrix_50_8 = 252'he4821045fa6784c0a499c22ad8697ffb20c43fe7abf2c1a844f8f8f9e3cc82d;
  assign mdsMatrix_51_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_51_1 = 253'h19199e443f564d1628b90e262a0c3dc6ea48ba435cc32b742bf02b53c8c700ef;
  assign mdsMatrix_51_2 = 255'h47d5b70845b435ea2ce4061441a1951396264526d3fca4e7b4a06fc33c80d9f8;
  assign mdsMatrix_51_3 = 254'h3e2c00494b673d9cb72c7ed47f5682014ced50236c51186193956916eb34b3b3;
  assign mdsMatrix_51_4 = 254'h34f97a52b8a7cc2157a2d6246a348502f39adb3eac33cb11265355d3e49c8356;
  assign mdsMatrix_51_5 = 253'h16f120d0fd9d217b1906f012851a3890aa5eb00761cc1542dbdbef08225514a4;
  assign mdsMatrix_51_6 = 255'h68be7d4c2805990ff7a838043424f9ba82a5efc1757993a1ee66df2f9ba745c5;
  assign mdsMatrix_51_7 = 255'h4a59bdc54a72b717a3ce99a87c27a6a7b5cffaf74998b37ede740b72e2798de3;
  assign mdsMatrix_51_8 = 255'h54e3e276dc63ccc4c1bce82b016b1f0c31f6a4a36ee4641cac7e948764283ead;
  assign mdsMatrix_52_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_52_1 = 255'h738644660b4e9b827752bc3d18fb698f2f86db6bb178c7f2ee95f559c069a78c;
  assign mdsMatrix_52_2 = 255'h42a7f6473657baa855520e5b0764a445327c4e28965efe5feb27346ff71d5eae;
  assign mdsMatrix_52_3 = 255'h65854fea633300572677a1bfdc231c1662e0ce05badc33a8f9698f54682c507d;
  assign mdsMatrix_52_4 = 254'h280349d42b5733d58cf833f47ae197331b47cd82232aff6937c8a4da97e6af25;
  assign mdsMatrix_52_5 = 255'h47c095c38e443c5e59949916c89826ddba3b3eca61ee914fe056af4b9fed5800;
  assign mdsMatrix_52_6 = 255'h409b4c754b90fc555b1fb1799fb892acc778b66794117339106d80b0bae99a78;
  assign mdsMatrix_52_7 = 255'h5782ee4504d51a09fc7f0bfc8b6473558c939dfd51a28dc5c7ead90a3610a393;
  assign mdsMatrix_52_8 = 253'h157ccf020fd0efa87519f2e8e0d8a1ac19ca1f9bd5f41adbda70c4c0627ddcad;
  assign mdsMatrix_53_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_53_1 = 254'h2de240fed108777af522ec355bae35f73097d185d8c759c558e4ee5416f426ca;
  assign mdsMatrix_53_2 = 253'h1017c2e25e2020f2da6f8f5dcc12f989860c2c28ec5cdf63fe21a34013acf370;
  assign mdsMatrix_53_3 = 255'h66dc261537fb9da49530334ecddb0a98ebbfa359926e5d9f6f3a4ebfd661f5ec;
  assign mdsMatrix_53_4 = 254'h2a598982cd29e52cb67867dca4125c20f863f99002656895e609616b45daa5d1;
  assign mdsMatrix_53_5 = 255'h5e04f006b21a8176e70000b39fde8ac66961e9395ea697b1c2e926722ea66fd7;
  assign mdsMatrix_53_6 = 254'h2b4579f433f0c92adf0af838f2902de6bcd133ecc2cd1e77154cc576ea46cb1e;
  assign mdsMatrix_53_7 = 254'h2aece527247818f3b0988bd244879428f13972a4eb17ecf5d6cb60c5f26fdd94;
  assign mdsMatrix_53_8 = 254'h2fbe3e41456527cd6c87fd448034fc6a6ebd2e2e5d79167ea6e6d0f3161ee927;
  assign mdsMatrix_54_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_54_1 = 253'h1a5ec0c84bf6c6403fb163c68b65d429ec80545153e85bd4bb9f1f81d1635bb4;
  assign mdsMatrix_54_2 = 255'h71ab0f88c4b5cf7e315805a26934f35cb7b6c7f5ddc7b072b4572d067198c426;
  assign mdsMatrix_54_3 = 255'h61e9a15fdbada59ed01895b171a05cc3306ffaa99a8f20bef22483c6c2569bf7;
  assign mdsMatrix_54_4 = 255'h69a08925816b2150762b3a2ba8f10ef92b12555c4d528d448ae919ae5a050da8;
  assign mdsMatrix_54_5 = 254'h21bc8468d55088b032d5ce33afb02ff1510a5a3d5fc02982adfa24b4dfd20caa;
  assign mdsMatrix_54_6 = 255'h4ac42147668103a4c031097d12dbc78e0e80d56abc0e5a1708f29f9ff4694184;
  assign mdsMatrix_54_7 = 253'h15dff9aada990b1a4a8819dd283627387605f52314bdeb49ff898f335fca1ff4;
  assign mdsMatrix_54_8 = 254'h3ed22826809e02fcb57f39053b5252cdea64df435606f1962d2a8377b855c9e2;
  assign mdsMatrix_55_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_55_1 = 252'hdf436eb17ae2a9b34569e6694200a7d4620a89f5b05a705aaaaaaaaa4fa4fa5;
  assign mdsMatrix_55_2 = 252'hd43617107703d62ad27b6d64b6715ea2f16e2859bc00cf4bc39293cd00a044d;
  assign mdsMatrix_55_3 = 255'h6346e1847f6c7c34119b8383de861dea1a65a6d87e958cb928261b7d1e9a96c8;
  assign mdsMatrix_55_4 = 255'h4cc1fcbd7729da5453b911245684982a3474c974e6e8a788fd0e83bcc7f30107;
  assign mdsMatrix_55_5 = 255'h4340b572ea97fe04723092792502007c6713b231c0b4bd7a2f83f7055d7743fb;
  assign mdsMatrix_55_6 = 255'h442d9b0cbc7d1ad713339a54a8eae39474946c1da1151942f9382c7588c18081;
  assign mdsMatrix_55_7 = 255'h463db9682b9ecd9aa79f744954c05dbcb50b2f56a27373bf67e70189384455c4;
  assign mdsMatrix_55_8 = 255'h6b3509dd57339338bf29f4140289fac58969d8ccbf626c912e1d548ae0be80f5;
  assign mdsMatrix_56_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_56_1 = 250'h26a11bc2ae0808b28f46e64cadfa19888da1265cccd20cd0000000033333333;
  assign mdsMatrix_56_2 = 254'h2c59c154f04b2e0d209627474791ca2f8396d8008ba29c5ce8ba2e8b745d1746;
  assign mdsMatrix_56_3 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_56_4 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_56_5 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_56_6 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_56_7 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_56_8 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign tempAddrVec_5 = io_addr_regNext_5;
  assign tempAddrVec_6 = io_addr_regNext_6;
  assign tempAddrVec_7 = io_addr_regNext_7;
  assign tempAddrVec_8 = io_addr_regNext_8;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  assign io_data_5 = _zz_mdsMem_5_port0;
  assign io_data_6 = _zz_mdsMem_6_port0;
  assign io_data_7 = _zz_mdsMem_7_port0;
  assign io_data_8 = _zz_mdsMem_8_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
    io_addr_regNext_5 <= io_addr;
    io_addr_regNext_6 <= io_addr;
    io_addr_regNext_7 <= io_addr;
    io_addr_regNext_8 <= io_addr;
  end


endmodule

module MatrixConstantMem_9 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  input      [5:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  reg        [254:0]  _zz_mdsMem_5_port0;
  reg        [254:0]  _zz_mdsMem_6_port0;
  reg        [254:0]  _zz_mdsMem_7_port0;
  reg        [254:0]  _zz_mdsMem_8_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire                _zz_mdsMem_5_port;
  wire                _zz_io_data_5;
  wire                _zz_mdsMem_6_port;
  wire                _zz_io_data_6;
  wire                _zz_mdsMem_7_port;
  wire                _zz_io_data_7;
  wire                _zz_mdsMem_8_port;
  wire                _zz_io_data_8;
  wire       [250:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [253:0]  mdsMatrix_0_2;
  wire       [250:0]  mdsMatrix_0_3;
  wire       [254:0]  mdsMatrix_0_4;
  wire       [250:0]  mdsMatrix_0_5;
  wire       [252:0]  mdsMatrix_0_6;
  wire       [254:0]  mdsMatrix_0_7;
  wire       [254:0]  mdsMatrix_0_8;
  wire       [250:0]  mdsMatrix_1_0;
  wire       [253:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [253:0]  mdsMatrix_1_3;
  wire       [253:0]  mdsMatrix_1_4;
  wire       [253:0]  mdsMatrix_1_5;
  wire       [254:0]  mdsMatrix_1_6;
  wire       [253:0]  mdsMatrix_1_7;
  wire       [251:0]  mdsMatrix_1_8;
  wire       [250:0]  mdsMatrix_2_0;
  wire       [253:0]  mdsMatrix_2_1;
  wire       [253:0]  mdsMatrix_2_2;
  wire       [254:0]  mdsMatrix_2_3;
  wire       [254:0]  mdsMatrix_2_4;
  wire       [252:0]  mdsMatrix_2_5;
  wire       [254:0]  mdsMatrix_2_6;
  wire       [253:0]  mdsMatrix_2_7;
  wire       [250:0]  mdsMatrix_2_8;
  wire       [250:0]  mdsMatrix_3_0;
  wire       [243:0]  mdsMatrix_3_1;
  wire       [254:0]  mdsMatrix_3_2;
  wire       [251:0]  mdsMatrix_3_3;
  wire       [252:0]  mdsMatrix_3_4;
  wire       [254:0]  mdsMatrix_3_5;
  wire       [252:0]  mdsMatrix_3_6;
  wire       [250:0]  mdsMatrix_3_7;
  wire       [254:0]  mdsMatrix_3_8;
  wire       [250:0]  mdsMatrix_4_0;
  wire       [254:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [253:0]  mdsMatrix_4_3;
  wire       [253:0]  mdsMatrix_4_4;
  wire       [254:0]  mdsMatrix_4_5;
  wire       [253:0]  mdsMatrix_4_6;
  wire       [254:0]  mdsMatrix_4_7;
  wire       [253:0]  mdsMatrix_4_8;
  wire       [250:0]  mdsMatrix_5_0;
  wire       [252:0]  mdsMatrix_5_1;
  wire       [252:0]  mdsMatrix_5_2;
  wire       [254:0]  mdsMatrix_5_3;
  wire       [253:0]  mdsMatrix_5_4;
  wire       [252:0]  mdsMatrix_5_5;
  wire       [253:0]  mdsMatrix_5_6;
  wire       [253:0]  mdsMatrix_5_7;
  wire       [254:0]  mdsMatrix_5_8;
  wire       [250:0]  mdsMatrix_6_0;
  wire       [253:0]  mdsMatrix_6_1;
  wire       [249:0]  mdsMatrix_6_2;
  wire       [252:0]  mdsMatrix_6_3;
  wire       [251:0]  mdsMatrix_6_4;
  wire       [254:0]  mdsMatrix_6_5;
  wire       [254:0]  mdsMatrix_6_6;
  wire       [252:0]  mdsMatrix_6_7;
  wire       [254:0]  mdsMatrix_6_8;
  wire       [250:0]  mdsMatrix_7_0;
  wire       [254:0]  mdsMatrix_7_1;
  wire       [254:0]  mdsMatrix_7_2;
  wire       [252:0]  mdsMatrix_7_3;
  wire       [250:0]  mdsMatrix_7_4;
  wire       [253:0]  mdsMatrix_7_5;
  wire       [252:0]  mdsMatrix_7_6;
  wire       [253:0]  mdsMatrix_7_7;
  wire       [254:0]  mdsMatrix_7_8;
  wire       [250:0]  mdsMatrix_8_0;
  wire       [253:0]  mdsMatrix_8_1;
  wire       [251:0]  mdsMatrix_8_2;
  wire       [254:0]  mdsMatrix_8_3;
  wire       [252:0]  mdsMatrix_8_4;
  wire       [254:0]  mdsMatrix_8_5;
  wire       [252:0]  mdsMatrix_8_6;
  wire       [253:0]  mdsMatrix_8_7;
  wire       [254:0]  mdsMatrix_8_8;
  wire       [250:0]  mdsMatrix_9_0;
  wire       [251:0]  mdsMatrix_9_1;
  wire       [254:0]  mdsMatrix_9_2;
  wire       [252:0]  mdsMatrix_9_3;
  wire       [251:0]  mdsMatrix_9_4;
  wire       [253:0]  mdsMatrix_9_5;
  wire       [253:0]  mdsMatrix_9_6;
  wire       [253:0]  mdsMatrix_9_7;
  wire       [252:0]  mdsMatrix_9_8;
  wire       [250:0]  mdsMatrix_10_0;
  wire       [254:0]  mdsMatrix_10_1;
  wire       [254:0]  mdsMatrix_10_2;
  wire       [253:0]  mdsMatrix_10_3;
  wire       [252:0]  mdsMatrix_10_4;
  wire       [253:0]  mdsMatrix_10_5;
  wire       [253:0]  mdsMatrix_10_6;
  wire       [251:0]  mdsMatrix_10_7;
  wire       [253:0]  mdsMatrix_10_8;
  wire       [250:0]  mdsMatrix_11_0;
  wire       [253:0]  mdsMatrix_11_1;
  wire       [254:0]  mdsMatrix_11_2;
  wire       [254:0]  mdsMatrix_11_3;
  wire       [254:0]  mdsMatrix_11_4;
  wire       [252:0]  mdsMatrix_11_5;
  wire       [254:0]  mdsMatrix_11_6;
  wire       [254:0]  mdsMatrix_11_7;
  wire       [254:0]  mdsMatrix_11_8;
  wire       [250:0]  mdsMatrix_12_0;
  wire       [253:0]  mdsMatrix_12_1;
  wire       [251:0]  mdsMatrix_12_2;
  wire       [242:0]  mdsMatrix_12_3;
  wire       [251:0]  mdsMatrix_12_4;
  wire       [253:0]  mdsMatrix_12_5;
  wire       [254:0]  mdsMatrix_12_6;
  wire       [252:0]  mdsMatrix_12_7;
  wire       [254:0]  mdsMatrix_12_8;
  wire       [250:0]  mdsMatrix_13_0;
  wire       [250:0]  mdsMatrix_13_1;
  wire       [253:0]  mdsMatrix_13_2;
  wire       [250:0]  mdsMatrix_13_3;
  wire       [250:0]  mdsMatrix_13_4;
  wire       [251:0]  mdsMatrix_13_5;
  wire       [254:0]  mdsMatrix_13_6;
  wire       [253:0]  mdsMatrix_13_7;
  wire       [253:0]  mdsMatrix_13_8;
  wire       [250:0]  mdsMatrix_14_0;
  wire       [254:0]  mdsMatrix_14_1;
  wire       [254:0]  mdsMatrix_14_2;
  wire       [254:0]  mdsMatrix_14_3;
  wire       [254:0]  mdsMatrix_14_4;
  wire       [254:0]  mdsMatrix_14_5;
  wire       [253:0]  mdsMatrix_14_6;
  wire       [254:0]  mdsMatrix_14_7;
  wire       [253:0]  mdsMatrix_14_8;
  wire       [250:0]  mdsMatrix_15_0;
  wire       [254:0]  mdsMatrix_15_1;
  wire       [254:0]  mdsMatrix_15_2;
  wire       [254:0]  mdsMatrix_15_3;
  wire       [253:0]  mdsMatrix_15_4;
  wire       [253:0]  mdsMatrix_15_5;
  wire       [252:0]  mdsMatrix_15_6;
  wire       [254:0]  mdsMatrix_15_7;
  wire       [254:0]  mdsMatrix_15_8;
  wire       [250:0]  mdsMatrix_16_0;
  wire       [251:0]  mdsMatrix_16_1;
  wire       [253:0]  mdsMatrix_16_2;
  wire       [252:0]  mdsMatrix_16_3;
  wire       [253:0]  mdsMatrix_16_4;
  wire       [254:0]  mdsMatrix_16_5;
  wire       [254:0]  mdsMatrix_16_6;
  wire       [252:0]  mdsMatrix_16_7;
  wire       [254:0]  mdsMatrix_16_8;
  wire       [250:0]  mdsMatrix_17_0;
  wire       [254:0]  mdsMatrix_17_1;
  wire       [253:0]  mdsMatrix_17_2;
  wire       [254:0]  mdsMatrix_17_3;
  wire       [254:0]  mdsMatrix_17_4;
  wire       [253:0]  mdsMatrix_17_5;
  wire       [254:0]  mdsMatrix_17_6;
  wire       [254:0]  mdsMatrix_17_7;
  wire       [254:0]  mdsMatrix_17_8;
  wire       [250:0]  mdsMatrix_18_0;
  wire       [252:0]  mdsMatrix_18_1;
  wire       [253:0]  mdsMatrix_18_2;
  wire       [252:0]  mdsMatrix_18_3;
  wire       [254:0]  mdsMatrix_18_4;
  wire       [254:0]  mdsMatrix_18_5;
  wire       [250:0]  mdsMatrix_18_6;
  wire       [253:0]  mdsMatrix_18_7;
  wire       [253:0]  mdsMatrix_18_8;
  wire       [250:0]  mdsMatrix_19_0;
  wire       [254:0]  mdsMatrix_19_1;
  wire       [251:0]  mdsMatrix_19_2;
  wire       [253:0]  mdsMatrix_19_3;
  wire       [253:0]  mdsMatrix_19_4;
  wire       [253:0]  mdsMatrix_19_5;
  wire       [254:0]  mdsMatrix_19_6;
  wire       [254:0]  mdsMatrix_19_7;
  wire       [254:0]  mdsMatrix_19_8;
  wire       [250:0]  mdsMatrix_20_0;
  wire       [254:0]  mdsMatrix_20_1;
  wire       [254:0]  mdsMatrix_20_2;
  wire       [253:0]  mdsMatrix_20_3;
  wire       [254:0]  mdsMatrix_20_4;
  wire       [254:0]  mdsMatrix_20_5;
  wire       [251:0]  mdsMatrix_20_6;
  wire       [252:0]  mdsMatrix_20_7;
  wire       [251:0]  mdsMatrix_20_8;
  wire       [250:0]  mdsMatrix_21_0;
  wire       [254:0]  mdsMatrix_21_1;
  wire       [252:0]  mdsMatrix_21_2;
  wire       [253:0]  mdsMatrix_21_3;
  wire       [252:0]  mdsMatrix_21_4;
  wire       [253:0]  mdsMatrix_21_5;
  wire       [254:0]  mdsMatrix_21_6;
  wire       [254:0]  mdsMatrix_21_7;
  wire       [253:0]  mdsMatrix_21_8;
  wire       [250:0]  mdsMatrix_22_0;
  wire       [253:0]  mdsMatrix_22_1;
  wire       [251:0]  mdsMatrix_22_2;
  wire       [254:0]  mdsMatrix_22_3;
  wire       [252:0]  mdsMatrix_22_4;
  wire       [254:0]  mdsMatrix_22_5;
  wire       [252:0]  mdsMatrix_22_6;
  wire       [253:0]  mdsMatrix_22_7;
  wire       [254:0]  mdsMatrix_22_8;
  wire       [250:0]  mdsMatrix_23_0;
  wire       [253:0]  mdsMatrix_23_1;
  wire       [254:0]  mdsMatrix_23_2;
  wire       [253:0]  mdsMatrix_23_3;
  wire       [254:0]  mdsMatrix_23_4;
  wire       [253:0]  mdsMatrix_23_5;
  wire       [254:0]  mdsMatrix_23_6;
  wire       [254:0]  mdsMatrix_23_7;
  wire       [252:0]  mdsMatrix_23_8;
  wire       [250:0]  mdsMatrix_24_0;
  wire       [251:0]  mdsMatrix_24_1;
  wire       [254:0]  mdsMatrix_24_2;
  wire       [253:0]  mdsMatrix_24_3;
  wire       [253:0]  mdsMatrix_24_4;
  wire       [252:0]  mdsMatrix_24_5;
  wire       [254:0]  mdsMatrix_24_6;
  wire       [253:0]  mdsMatrix_24_7;
  wire       [252:0]  mdsMatrix_24_8;
  wire       [250:0]  mdsMatrix_25_0;
  wire       [254:0]  mdsMatrix_25_1;
  wire       [250:0]  mdsMatrix_25_2;
  wire       [254:0]  mdsMatrix_25_3;
  wire       [250:0]  mdsMatrix_25_4;
  wire       [253:0]  mdsMatrix_25_5;
  wire       [254:0]  mdsMatrix_25_6;
  wire       [254:0]  mdsMatrix_25_7;
  wire       [253:0]  mdsMatrix_25_8;
  wire       [250:0]  mdsMatrix_26_0;
  wire       [253:0]  mdsMatrix_26_1;
  wire       [252:0]  mdsMatrix_26_2;
  wire       [250:0]  mdsMatrix_26_3;
  wire       [254:0]  mdsMatrix_26_4;
  wire       [254:0]  mdsMatrix_26_5;
  wire       [253:0]  mdsMatrix_26_6;
  wire       [253:0]  mdsMatrix_26_7;
  wire       [254:0]  mdsMatrix_26_8;
  wire       [250:0]  mdsMatrix_27_0;
  wire       [253:0]  mdsMatrix_27_1;
  wire       [254:0]  mdsMatrix_27_2;
  wire       [254:0]  mdsMatrix_27_3;
  wire       [254:0]  mdsMatrix_27_4;
  wire       [254:0]  mdsMatrix_27_5;
  wire       [254:0]  mdsMatrix_27_6;
  wire       [251:0]  mdsMatrix_27_7;
  wire       [249:0]  mdsMatrix_27_8;
  wire       [250:0]  mdsMatrix_28_0;
  wire       [254:0]  mdsMatrix_28_1;
  wire       [252:0]  mdsMatrix_28_2;
  wire       [251:0]  mdsMatrix_28_3;
  wire       [254:0]  mdsMatrix_28_4;
  wire       [254:0]  mdsMatrix_28_5;
  wire       [254:0]  mdsMatrix_28_6;
  wire       [253:0]  mdsMatrix_28_7;
  wire       [254:0]  mdsMatrix_28_8;
  wire       [250:0]  mdsMatrix_29_0;
  wire       [254:0]  mdsMatrix_29_1;
  wire       [253:0]  mdsMatrix_29_2;
  wire       [254:0]  mdsMatrix_29_3;
  wire       [254:0]  mdsMatrix_29_4;
  wire       [253:0]  mdsMatrix_29_5;
  wire       [253:0]  mdsMatrix_29_6;
  wire       [254:0]  mdsMatrix_29_7;
  wire       [253:0]  mdsMatrix_29_8;
  wire       [250:0]  mdsMatrix_30_0;
  wire       [253:0]  mdsMatrix_30_1;
  wire       [253:0]  mdsMatrix_30_2;
  wire       [252:0]  mdsMatrix_30_3;
  wire       [254:0]  mdsMatrix_30_4;
  wire       [254:0]  mdsMatrix_30_5;
  wire       [254:0]  mdsMatrix_30_6;
  wire       [253:0]  mdsMatrix_30_7;
  wire       [252:0]  mdsMatrix_30_8;
  wire       [250:0]  mdsMatrix_31_0;
  wire       [252:0]  mdsMatrix_31_1;
  wire       [253:0]  mdsMatrix_31_2;
  wire       [252:0]  mdsMatrix_31_3;
  wire       [254:0]  mdsMatrix_31_4;
  wire       [253:0]  mdsMatrix_31_5;
  wire       [254:0]  mdsMatrix_31_6;
  wire       [254:0]  mdsMatrix_31_7;
  wire       [253:0]  mdsMatrix_31_8;
  wire       [250:0]  mdsMatrix_32_0;
  wire       [253:0]  mdsMatrix_32_1;
  wire       [254:0]  mdsMatrix_32_2;
  wire       [254:0]  mdsMatrix_32_3;
  wire       [252:0]  mdsMatrix_32_4;
  wire       [253:0]  mdsMatrix_32_5;
  wire       [251:0]  mdsMatrix_32_6;
  wire       [254:0]  mdsMatrix_32_7;
  wire       [251:0]  mdsMatrix_32_8;
  wire       [250:0]  mdsMatrix_33_0;
  wire       [252:0]  mdsMatrix_33_1;
  wire       [254:0]  mdsMatrix_33_2;
  wire       [253:0]  mdsMatrix_33_3;
  wire       [254:0]  mdsMatrix_33_4;
  wire       [253:0]  mdsMatrix_33_5;
  wire       [252:0]  mdsMatrix_33_6;
  wire       [251:0]  mdsMatrix_33_7;
  wire       [254:0]  mdsMatrix_33_8;
  wire       [250:0]  mdsMatrix_34_0;
  wire       [254:0]  mdsMatrix_34_1;
  wire       [252:0]  mdsMatrix_34_2;
  wire       [250:0]  mdsMatrix_34_3;
  wire       [254:0]  mdsMatrix_34_4;
  wire       [254:0]  mdsMatrix_34_5;
  wire       [254:0]  mdsMatrix_34_6;
  wire       [254:0]  mdsMatrix_34_7;
  wire       [252:0]  mdsMatrix_34_8;
  wire       [250:0]  mdsMatrix_35_0;
  wire       [254:0]  mdsMatrix_35_1;
  wire       [254:0]  mdsMatrix_35_2;
  wire       [254:0]  mdsMatrix_35_3;
  wire       [254:0]  mdsMatrix_35_4;
  wire       [252:0]  mdsMatrix_35_5;
  wire       [254:0]  mdsMatrix_35_6;
  wire       [254:0]  mdsMatrix_35_7;
  wire       [252:0]  mdsMatrix_35_8;
  wire       [250:0]  mdsMatrix_36_0;
  wire       [252:0]  mdsMatrix_36_1;
  wire       [254:0]  mdsMatrix_36_2;
  wire       [254:0]  mdsMatrix_36_3;
  wire       [254:0]  mdsMatrix_36_4;
  wire       [254:0]  mdsMatrix_36_5;
  wire       [250:0]  mdsMatrix_36_6;
  wire       [253:0]  mdsMatrix_36_7;
  wire       [253:0]  mdsMatrix_36_8;
  wire       [250:0]  mdsMatrix_37_0;
  wire       [254:0]  mdsMatrix_37_1;
  wire       [254:0]  mdsMatrix_37_2;
  wire       [254:0]  mdsMatrix_37_3;
  wire       [254:0]  mdsMatrix_37_4;
  wire       [253:0]  mdsMatrix_37_5;
  wire       [254:0]  mdsMatrix_37_6;
  wire       [253:0]  mdsMatrix_37_7;
  wire       [254:0]  mdsMatrix_37_8;
  wire       [250:0]  mdsMatrix_38_0;
  wire       [254:0]  mdsMatrix_38_1;
  wire       [254:0]  mdsMatrix_38_2;
  wire       [254:0]  mdsMatrix_38_3;
  wire       [254:0]  mdsMatrix_38_4;
  wire       [249:0]  mdsMatrix_38_5;
  wire       [253:0]  mdsMatrix_38_6;
  wire       [254:0]  mdsMatrix_38_7;
  wire       [254:0]  mdsMatrix_38_8;
  wire       [250:0]  mdsMatrix_39_0;
  wire       [252:0]  mdsMatrix_39_1;
  wire       [254:0]  mdsMatrix_39_2;
  wire       [249:0]  mdsMatrix_39_3;
  wire       [254:0]  mdsMatrix_39_4;
  wire       [254:0]  mdsMatrix_39_5;
  wire       [253:0]  mdsMatrix_39_6;
  wire       [254:0]  mdsMatrix_39_7;
  wire       [254:0]  mdsMatrix_39_8;
  wire       [250:0]  mdsMatrix_40_0;
  wire       [253:0]  mdsMatrix_40_1;
  wire       [254:0]  mdsMatrix_40_2;
  wire       [253:0]  mdsMatrix_40_3;
  wire       [253:0]  mdsMatrix_40_4;
  wire       [254:0]  mdsMatrix_40_5;
  wire       [254:0]  mdsMatrix_40_6;
  wire       [254:0]  mdsMatrix_40_7;
  wire       [254:0]  mdsMatrix_40_8;
  wire       [250:0]  mdsMatrix_41_0;
  wire       [251:0]  mdsMatrix_41_1;
  wire       [253:0]  mdsMatrix_41_2;
  wire       [254:0]  mdsMatrix_41_3;
  wire       [253:0]  mdsMatrix_41_4;
  wire       [254:0]  mdsMatrix_41_5;
  wire       [252:0]  mdsMatrix_41_6;
  wire       [250:0]  mdsMatrix_41_7;
  wire       [253:0]  mdsMatrix_41_8;
  wire       [250:0]  mdsMatrix_42_0;
  wire       [252:0]  mdsMatrix_42_1;
  wire       [254:0]  mdsMatrix_42_2;
  wire       [254:0]  mdsMatrix_42_3;
  wire       [254:0]  mdsMatrix_42_4;
  wire       [252:0]  mdsMatrix_42_5;
  wire       [253:0]  mdsMatrix_42_6;
  wire       [253:0]  mdsMatrix_42_7;
  wire       [254:0]  mdsMatrix_42_8;
  wire       [250:0]  mdsMatrix_43_0;
  wire       [254:0]  mdsMatrix_43_1;
  wire       [251:0]  mdsMatrix_43_2;
  wire       [253:0]  mdsMatrix_43_3;
  wire       [253:0]  mdsMatrix_43_4;
  wire       [252:0]  mdsMatrix_43_5;
  wire       [253:0]  mdsMatrix_43_6;
  wire       [253:0]  mdsMatrix_43_7;
  wire       [251:0]  mdsMatrix_43_8;
  wire       [250:0]  mdsMatrix_44_0;
  wire       [251:0]  mdsMatrix_44_1;
  wire       [253:0]  mdsMatrix_44_2;
  wire       [252:0]  mdsMatrix_44_3;
  wire       [254:0]  mdsMatrix_44_4;
  wire       [253:0]  mdsMatrix_44_5;
  wire       [254:0]  mdsMatrix_44_6;
  wire       [254:0]  mdsMatrix_44_7;
  wire       [254:0]  mdsMatrix_44_8;
  wire       [250:0]  mdsMatrix_45_0;
  wire       [254:0]  mdsMatrix_45_1;
  wire       [254:0]  mdsMatrix_45_2;
  wire       [253:0]  mdsMatrix_45_3;
  wire       [249:0]  mdsMatrix_45_4;
  wire       [250:0]  mdsMatrix_45_5;
  wire       [252:0]  mdsMatrix_45_6;
  wire       [254:0]  mdsMatrix_45_7;
  wire       [254:0]  mdsMatrix_45_8;
  wire       [250:0]  mdsMatrix_46_0;
  wire       [253:0]  mdsMatrix_46_1;
  wire       [251:0]  mdsMatrix_46_2;
  wire       [254:0]  mdsMatrix_46_3;
  wire       [253:0]  mdsMatrix_46_4;
  wire       [254:0]  mdsMatrix_46_5;
  wire       [254:0]  mdsMatrix_46_6;
  wire       [254:0]  mdsMatrix_46_7;
  wire       [254:0]  mdsMatrix_46_8;
  wire       [250:0]  mdsMatrix_47_0;
  wire       [253:0]  mdsMatrix_47_1;
  wire       [251:0]  mdsMatrix_47_2;
  wire       [253:0]  mdsMatrix_47_3;
  wire       [252:0]  mdsMatrix_47_4;
  wire       [253:0]  mdsMatrix_47_5;
  wire       [254:0]  mdsMatrix_47_6;
  wire       [250:0]  mdsMatrix_47_7;
  wire       [253:0]  mdsMatrix_47_8;
  wire       [250:0]  mdsMatrix_48_0;
  wire       [254:0]  mdsMatrix_48_1;
  wire       [254:0]  mdsMatrix_48_2;
  wire       [254:0]  mdsMatrix_48_3;
  wire       [253:0]  mdsMatrix_48_4;
  wire       [254:0]  mdsMatrix_48_5;
  wire       [250:0]  mdsMatrix_48_6;
  wire       [253:0]  mdsMatrix_48_7;
  wire       [254:0]  mdsMatrix_48_8;
  wire       [250:0]  mdsMatrix_49_0;
  wire       [252:0]  mdsMatrix_49_1;
  wire       [252:0]  mdsMatrix_49_2;
  wire       [254:0]  mdsMatrix_49_3;
  wire       [254:0]  mdsMatrix_49_4;
  wire       [251:0]  mdsMatrix_49_5;
  wire       [253:0]  mdsMatrix_49_6;
  wire       [254:0]  mdsMatrix_49_7;
  wire       [254:0]  mdsMatrix_49_8;
  wire       [250:0]  mdsMatrix_50_0;
  wire       [253:0]  mdsMatrix_50_1;
  wire       [252:0]  mdsMatrix_50_2;
  wire       [254:0]  mdsMatrix_50_3;
  wire       [254:0]  mdsMatrix_50_4;
  wire       [253:0]  mdsMatrix_50_5;
  wire       [253:0]  mdsMatrix_50_6;
  wire       [251:0]  mdsMatrix_50_7;
  wire       [251:0]  mdsMatrix_50_8;
  wire       [250:0]  mdsMatrix_51_0;
  wire       [251:0]  mdsMatrix_51_1;
  wire       [251:0]  mdsMatrix_51_2;
  wire       [250:0]  mdsMatrix_51_3;
  wire       [253:0]  mdsMatrix_51_4;
  wire       [254:0]  mdsMatrix_51_5;
  wire       [254:0]  mdsMatrix_51_6;
  wire       [252:0]  mdsMatrix_51_7;
  wire       [252:0]  mdsMatrix_51_8;
  wire       [250:0]  mdsMatrix_52_0;
  wire       [253:0]  mdsMatrix_52_1;
  wire       [253:0]  mdsMatrix_52_2;
  wire       [254:0]  mdsMatrix_52_3;
  wire       [253:0]  mdsMatrix_52_4;
  wire       [253:0]  mdsMatrix_52_5;
  wire       [251:0]  mdsMatrix_52_6;
  wire       [254:0]  mdsMatrix_52_7;
  wire       [253:0]  mdsMatrix_52_8;
  wire       [250:0]  mdsMatrix_53_0;
  wire       [251:0]  mdsMatrix_53_1;
  wire       [254:0]  mdsMatrix_53_2;
  wire       [253:0]  mdsMatrix_53_3;
  wire       [253:0]  mdsMatrix_53_4;
  wire       [251:0]  mdsMatrix_53_5;
  wire       [254:0]  mdsMatrix_53_6;
  wire       [254:0]  mdsMatrix_53_7;
  wire       [252:0]  mdsMatrix_53_8;
  wire       [250:0]  mdsMatrix_54_0;
  wire       [254:0]  mdsMatrix_54_1;
  wire       [254:0]  mdsMatrix_54_2;
  wire       [253:0]  mdsMatrix_54_3;
  wire       [254:0]  mdsMatrix_54_4;
  wire       [254:0]  mdsMatrix_54_5;
  wire       [252:0]  mdsMatrix_54_6;
  wire       [253:0]  mdsMatrix_54_7;
  wire       [251:0]  mdsMatrix_54_8;
  wire       [250:0]  mdsMatrix_55_0;
  wire       [254:0]  mdsMatrix_55_1;
  wire       [254:0]  mdsMatrix_55_2;
  wire       [253:0]  mdsMatrix_55_3;
  wire       [254:0]  mdsMatrix_55_4;
  wire       [250:0]  mdsMatrix_55_5;
  wire       [253:0]  mdsMatrix_55_6;
  wire       [254:0]  mdsMatrix_55_7;
  wire       [254:0]  mdsMatrix_55_8;
  wire       [5:0]    tempAddrVec_0;
  wire       [5:0]    tempAddrVec_1;
  wire       [5:0]    tempAddrVec_2;
  wire       [5:0]    tempAddrVec_3;
  wire       [5:0]    tempAddrVec_4;
  wire       [5:0]    tempAddrVec_5;
  wire       [5:0]    tempAddrVec_6;
  wire       [5:0]    tempAddrVec_7;
  wire       [5:0]    tempAddrVec_8;
  reg        [5:0]    io_addr_regNext;
  reg        [5:0]    io_addr_regNext_1;
  reg        [5:0]    io_addr_regNext_2;
  reg        [5:0]    io_addr_regNext_3;
  reg        [5:0]    io_addr_regNext_4;
  reg        [5:0]    io_addr_regNext_5;
  reg        [5:0]    io_addr_regNext_6;
  reg        [5:0]    io_addr_regNext_7;
  reg        [5:0]    io_addr_regNext_8;
  reg [254:0] mdsMem_0 [0:55];
  reg [254:0] mdsMem_1 [0:55];
  reg [254:0] mdsMem_2 [0:55];
  reg [254:0] mdsMem_3 [0:55];
  reg [254:0] mdsMem_4 [0:55];
  reg [254:0] mdsMem_5 [0:55];
  reg [254:0] mdsMem_6 [0:55];
  reg [254:0] mdsMem_7 [0:55];
  reg [254:0] mdsMem_8 [0:55];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  assign _zz_io_data_5 = 1'b1;
  assign _zz_io_data_6 = 1'b1;
  assign _zz_io_data_7 = 1'b1;
  assign _zz_io_data_8 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_23_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_23_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_23_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_23_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_23_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_23_mdsMem_5.bin",mdsMem_5);
  end
  always @(posedge clk) begin
    if(_zz_io_data_5) begin
      _zz_mdsMem_5_port0 <= mdsMem_5[tempAddrVec_5];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_23_mdsMem_6.bin",mdsMem_6);
  end
  always @(posedge clk) begin
    if(_zz_io_data_6) begin
      _zz_mdsMem_6_port0 <= mdsMem_6[tempAddrVec_6];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_23_mdsMem_7.bin",mdsMem_7);
  end
  always @(posedge clk) begin
    if(_zz_io_data_7) begin
      _zz_mdsMem_7_port0 <= mdsMem_7[tempAddrVec_7];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_23_mdsMem_8.bin",mdsMem_8);
  end
  always @(posedge clk) begin
    if(_zz_io_data_8) begin
      _zz_mdsMem_8_port0 <= mdsMem_8[tempAddrVec_8];
    end
  end

  assign mdsMatrix_0_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_0_1 = 255'h59f4fe1a17ec4ae7d1e34cc44c0d2007363fb23be4011de71f42e26f5cb19cc3;
  assign mdsMatrix_0_2 = 254'h3dbc31f0b557e434b17ec0c982dad58b85cd2df59f157ae99787462613220213;
  assign mdsMatrix_0_3 = 251'h45148a86ae553e26c3c9b5a4863c8a0568644136b24fc4890da028c7d7475c7;
  assign mdsMatrix_0_4 = 255'h498a8d4d62df169fe32dd32a7c8e30a4c076035058417e97b62cff3595aa5f93;
  assign mdsMatrix_0_5 = 251'h79f45ba66a03cc54768db87d6c2cc6bd4036676ba2f235a43962d041e587418;
  assign mdsMatrix_0_6 = 253'h18f1bf1ec04ad5a0ba4f75435de6fd95eeb86a7d310a58c1e3a87f755bc2b049;
  assign mdsMatrix_0_7 = 255'h42926696988d6a0221e5cbf2a1d430c5dfd83639be854c2fea6e0e3af008d77e;
  assign mdsMatrix_0_8 = 255'h4423453d163b940cf39cb29c1a84e821f1c3c6dd8955a9349059f783e4828624;
  assign mdsMatrix_1_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_1_1 = 254'h36881382839aa4cb6bb10a63971d68b8b77ccfedef598466822f7001d6634439;
  assign mdsMatrix_1_2 = 255'h586a13a470f5966adebd693d041b6169980f5005d43febfe6ae03dae387a4357;
  assign mdsMatrix_1_3 = 254'h24ca96cd9a66dc8308019a68101a59e311d935296fdddb12e1ffc06502e91cff;
  assign mdsMatrix_1_4 = 254'h3bce8276e15beb9c496c8f1b1cfb535fd499752376311297ce2ec437d6a5f671;
  assign mdsMatrix_1_5 = 254'h38ec1e8b0b3fa8e6a3271ad72fa8dc8245f12963c36cc6de1c0143cafe7b7059;
  assign mdsMatrix_1_6 = 255'h5cecb61bd21c25d437fecca36feddf6649fe87cb213b87f234dae05546eb5ebd;
  assign mdsMatrix_1_7 = 254'h2a96fe47bf1588d8ba3a9d0691cf64a18a72283052ed91448f42cfe0714632b2;
  assign mdsMatrix_1_8 = 252'hafb437c121d317c91d57aa84facb3a7be42dfd20803c266ae8c3c0137ff9b91;
  assign mdsMatrix_2_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_2_1 = 254'h32b0d04a7ce17d0497f95e592020036eb449c09b31f66fed24b0dc937a982a05;
  assign mdsMatrix_2_2 = 254'h39d0fa03aad43aaf95df985bc0049bb1b8922066f396c934fae64cfbb8b505f1;
  assign mdsMatrix_2_3 = 255'h522b9b823758b065dec2c17c5adea51a1fba7c61f811226284950c4fc19b8386;
  assign mdsMatrix_2_4 = 255'h50b169377a3f461dc901a7b554515ae7a6e58cd3941cfe19fd2263c2b5c97c3f;
  assign mdsMatrix_2_5 = 253'h1c04102cc202d989c2a8e9d4578861960a9c78f15118d4714af6e118e01dd351;
  assign mdsMatrix_2_6 = 255'h4285a04eb3edf30996e96ad0797ff69e095ca977408cb96bda92d31b9cc3504f;
  assign mdsMatrix_2_7 = 254'h3c46c34bd9757286dced0a46d42c50fffdf0ddeb76f6834272b4b7ac4323d804;
  assign mdsMatrix_2_8 = 251'h4362f93c5c980386cc49fbd335d82c278f02e44206b3b7c87f7a762bd56321f;
  assign mdsMatrix_3_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_3_1 = 244'hae5d86b3e8c2587a36a533074906b61443f6a703aefd4ca3a35dd2c6f584b;
  assign mdsMatrix_3_2 = 255'h5f8017198671956866141a55cf80dc8a26583689519fd817b638609a59b92dbf;
  assign mdsMatrix_3_3 = 252'hebc660e1c7df8753d6f6d417653bf3eb33f854b324b0e0160966ffd3335d1a3;
  assign mdsMatrix_3_4 = 253'h106969d0dbfed1f00e66b482ff52ec41261635c6e21a91817eeae1bbce1c00e4;
  assign mdsMatrix_3_5 = 255'h4bb2b70a69b5a30b1fae6a5749accb60be9b9f6e8776983b131096580e01747b;
  assign mdsMatrix_3_6 = 253'h1ba34a2f1a54898a3d088414db02620b383d74ebd060e35ce50f39e586f9aa8e;
  assign mdsMatrix_3_7 = 251'h757186627bd0d5412008c1f4b66b7f72745692efd4e4a5605453980e9417b13;
  assign mdsMatrix_3_8 = 255'h4c7bdfc617c113d81d7bb386a8ff3b9c4e2d13391ef2606b9728386517b40c12;
  assign mdsMatrix_4_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_4_1 = 255'h5d5be91b6796f04aaecafef9de1e4eb27189f47106de6878006d65ad4763160a;
  assign mdsMatrix_4_2 = 255'h7121bc6a928ab40e9cb267f5d18f6c46e964c5a10fbafb51aff8495db6e8c9d2;
  assign mdsMatrix_4_3 = 254'h3d61c506afc95e0321179376b46c388628cc9472eba0697ad5c82cf32502164c;
  assign mdsMatrix_4_4 = 254'h30778817e3281186d7d7453ddde1dda0492f77657aef296c685b245b5be9a3ff;
  assign mdsMatrix_4_5 = 255'h45614c2165276cc94945826925641f1a874c6267bb0fd184b6fb293ffad7c83f;
  assign mdsMatrix_4_6 = 254'h2890f578562455393790eb6648f117c400ebc659ce3fc353c0786dcca5614136;
  assign mdsMatrix_4_7 = 255'h495e92332fc918e8ab84b6019e441603bdfd04f3c0777a428e2e3d1f757d99a5;
  assign mdsMatrix_4_8 = 254'h2f57cecb5789c12ba3fc31c10c91176657ba59d4a6a46b7479e3f438d8ab2231;
  assign mdsMatrix_5_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_5_1 = 253'h1364780eb22a3fd97c29de841b1ec6c6ab36ffd879314bca99906f4b62b22320;
  assign mdsMatrix_5_2 = 253'h13cc3bfaf3153dd8c07d1fd9513ce2ccffb3e6b51befc9a6c49f43dd8e6d30cb;
  assign mdsMatrix_5_3 = 255'h6c371cb9e71e9ae75baa62228c5a0713f121ab9ec11629312e79798f0de8033c;
  assign mdsMatrix_5_4 = 254'h245924ba3f3ac458c0c13022c3aa9ec7762653179e22590086974c2046910508;
  assign mdsMatrix_5_5 = 253'h1847c981ea0e998169a204312cfd8125406908aacedf0efa8f19a293db067f0a;
  assign mdsMatrix_5_6 = 254'h2fa035591efc2aae83e0acb6461b65e6dbd0c5c52e6e6e288cfdd92d40c1c466;
  assign mdsMatrix_5_7 = 254'h3015825daa03222ac425ddd1f2bd999d5d924225e877fe766e1ca0cee8907492;
  assign mdsMatrix_5_8 = 255'h7100b7704ba2c0f130a54dd59dec85214515c49b3b073fbd443574467e217e28;
  assign mdsMatrix_6_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_6_1 = 254'h208bfd4bfe0d65ced70128e280bdc8a7a4129ea61495f513abab0031409105ce;
  assign mdsMatrix_6_2 = 250'h34d697627ecbbcadce655c48e7642fefc2842039387621d937fa6d74e23c3f0;
  assign mdsMatrix_6_3 = 253'h1fa111c90854b08575ef3f1ec5260b29e2f296166aa7b6a3a5b982676310bc91;
  assign mdsMatrix_6_4 = 252'hc787f6fb5558170817c5e45f2f74f9c73f20cefbfdc21b9007e4f9c0f7b361a;
  assign mdsMatrix_6_5 = 255'h4681064107e4d93caf30ef387314d62ab593907d1885a9bbc3e3fee6a8260c17;
  assign mdsMatrix_6_6 = 255'h59beb5da440af348a2dafd02a12f2ca8aca320db10b3be1dc7f82251748d855d;
  assign mdsMatrix_6_7 = 253'h18feea0a6bcdf8952c7538ac28f465d5761fefebed680be78642520fde456125;
  assign mdsMatrix_6_8 = 255'h6c10ba8cc8acef7694823f1f74299aecfe7c97c5f1790398d63eee053c08f334;
  assign mdsMatrix_7_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_7_1 = 255'h5a822bb118ec49c7d2c3a22a0a396a3b708a1f1697690f609e0cc8db4ee74212;
  assign mdsMatrix_7_2 = 255'h71a288f20c2dc725cb8c32a3a73f3ebafd699be1e58a482420646b74151bbca4;
  assign mdsMatrix_7_3 = 253'h15a8ad4bd35734eb7c3716deca84bf72802b91e51e9a456be4ccc8e6709f3284;
  assign mdsMatrix_7_4 = 251'h623c4fd4e698d4059bdc23ed1f257b7162a98ab9933a817e101caa75ceac6f8;
  assign mdsMatrix_7_5 = 254'h3ffe7a6760eea6ba6cecc596d50a8b64ba77a477a5d4513c210b1dbcd00f11a7;
  assign mdsMatrix_7_6 = 253'h19575a22430c473e74ef8387b1d52a1619a9a8391bdbc871fa2532d87adfb913;
  assign mdsMatrix_7_7 = 254'h3edd53eb8973f4b58cb756c36db7275772ef6ba820c7eacd9fbdad9a0b334a8d;
  assign mdsMatrix_7_8 = 255'h6bd957b249b809d790832fbfade158d3c7999ae5fded72a2ab2db311d22da328;
  assign mdsMatrix_8_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_8_1 = 254'h27faa7ca9be2ac56008e72d532152b0bd03bebb5f3193c71e7fc4a5575175766;
  assign mdsMatrix_8_2 = 252'hafc586f99ec81efbf33b650c317fb3aeafd5900479c25693e90a78d604b2875;
  assign mdsMatrix_8_3 = 255'h69c09ef2a36fc8e7ee9f6040adfa53da7ab8665460e44560136769304c2fc4bc;
  assign mdsMatrix_8_4 = 253'h168c084ba746b3a25816e5641775f4d3f2ca4366cec4a2ba1dd54ca75db1ac2f;
  assign mdsMatrix_8_5 = 255'h61c018a589bc82ad2ba3a0ce7ef9d3dd9eb25d25ffb894f16144a861be91d416;
  assign mdsMatrix_8_6 = 253'h1996a753689323703b92207c454f29498fbc712cc4288420769a82fd64cef1e8;
  assign mdsMatrix_8_7 = 254'h33659ad0cd1cf4bc8fb8301ee7b8c381326215b7b4fa950e269895a341b42a44;
  assign mdsMatrix_8_8 = 255'h632f8ad9d2328477cc3fa7648b18477c9e6c60fb80b553a8c39f200bad2b2572;
  assign mdsMatrix_9_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_9_1 = 252'hb136b1ae68b242d8406fe9f7b70a0fb07440144544b76f109d6c9eb679478f5;
  assign mdsMatrix_9_2 = 255'h60c7dd2abbdd9167791a279b3a5930cef837037d11c3e73ea2f336a9741739a5;
  assign mdsMatrix_9_3 = 253'h16072c9d744647dac401dcacd8cb3c33640f42d2231fe1b4fd4f780fe4a2e3b7;
  assign mdsMatrix_9_4 = 252'hbb88601ad86f6a37ebfc64b02ff4484354aca6e30f661b2ff3208558e434a65;
  assign mdsMatrix_9_5 = 254'h35c50e14a84e06aa32cf726b84cfd8dc825c97bb7739335470b6109374c2905b;
  assign mdsMatrix_9_6 = 254'h332cb671ee8948e3424998992fe5b411c17be4eb933c1439121546cdbd898139;
  assign mdsMatrix_9_7 = 254'h262f593579a3099226bf968ff6084c8a90b3223bda135bdd0604923703f32ed5;
  assign mdsMatrix_9_8 = 253'h14eef303a0ffc2a36ec20c74dfa7dcab00e09084d2244ef16479c5e0c7836c43;
  assign mdsMatrix_10_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_10_1 = 255'h6672a5580153b847452f5b14453e8f0130dd3c7d66e541c300b34d288bddc18f;
  assign mdsMatrix_10_2 = 255'h493f6f31839e9ef19fb71309a277390f7558201c878d789e3901c34a22c7f361;
  assign mdsMatrix_10_3 = 254'h380e6dec0cd9fbe62939e2d2088ed0ad60c9b0f34ba75013013ddd218d22b30e;
  assign mdsMatrix_10_4 = 253'h1208e92d2777aa44081c058716cb1c1b8c46782d0cba691189836797f085c952;
  assign mdsMatrix_10_5 = 254'h376c40268dc1d16d3d881b346d92523f5b2b9e81e42f1360095ec9f7f91aefa0;
  assign mdsMatrix_10_6 = 254'h34fec200df3294132af007b13c82f1aed5ff5ce6c4ae4d5334464404dde153c7;
  assign mdsMatrix_10_7 = 252'hed80d1674ed6cdee97256631f35979b74db1885433f32b6cb3a4304fa7adc47;
  assign mdsMatrix_10_8 = 254'h2c512be860545d210080c01118f15db989f69ba73e2652ec65d2ff9362a5b755;
  assign mdsMatrix_11_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_11_1 = 254'h3a5e19f827468b10f9e0de2d083a71912cd2c8ad19b5f8d47363e0f6848f0501;
  assign mdsMatrix_11_2 = 255'h44adb2be41ecaaa8ba6cd1f52ea1e0d005a1f2191acf0b2ff337388decb43ad6;
  assign mdsMatrix_11_3 = 255'h55c0555d77f0ac87b718a1dc9396c361c77754cf81d10d11d9b9dbe4b9c4949d;
  assign mdsMatrix_11_4 = 255'h44ffc21566f9580e407385546d71c03e6112382e45e092e6bf3524ac37d454aa;
  assign mdsMatrix_11_5 = 253'h195c7f7862fda6e4ee9bb6fa712dd6746c4686d4bea40ca5dba20cdc533d5289;
  assign mdsMatrix_11_6 = 255'h49b7a816824d7b540a5b0827cec419cfc21e3927e7cc6bb8fc7a6ef6d8d6762b;
  assign mdsMatrix_11_7 = 255'h5c706674323e0c42012cbdfa83b8ca5a0f27aa5abcf6f620eeacf6b10a439234;
  assign mdsMatrix_11_8 = 255'h66faa98c7ef890e04c6b2c3bd346c2d0340514184a87ae63980ae7a8521b2ffd;
  assign mdsMatrix_12_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_12_1 = 254'h271c257494cf510dbc4a708b658a9f4080ceaae7cb3d7a62e19b433609db7851;
  assign mdsMatrix_12_2 = 252'hbee15d195b6bae4148ac095f52544209416ef654a698a433c797368be09bbc8;
  assign mdsMatrix_12_3 = 243'h4a7a1f6e46a1f51b474058d7bb92ab49664b3a8435ec6725e88b5db33000f;
  assign mdsMatrix_12_4 = 252'ha84010a3362f4543ab8e90a8be9790d0b53f081150a71e24738e5063e671235;
  assign mdsMatrix_12_5 = 254'h3af0402eb27555bf464883f701fb4409e401eb22a27906913e803fa43d3fac8f;
  assign mdsMatrix_12_6 = 255'h41202e6f1f68ebe711a2409b696438da5464afc8d3b96298a08ef9dac6135339;
  assign mdsMatrix_12_7 = 253'h1a0ff7653ad19756ac22107fc1b6e5810428594b5e41b8591637ac6e327939cd;
  assign mdsMatrix_12_8 = 255'h412753981815afce05cbd319dfe619373eb95b64d642827bd74d516078cf3d75;
  assign mdsMatrix_13_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_13_1 = 251'h632c1e2ff1118466e95d874274dc0af3863faa4b02f8e5c352087285881f448;
  assign mdsMatrix_13_2 = 254'h350e045b1c71eb9d71441095ea98385105f460e1399b68adbf64c0e1143ff940;
  assign mdsMatrix_13_3 = 251'h6ebc528d582f91f8a17d2c89ae7f9181e729a78845c5ce45740fb91176e95ec;
  assign mdsMatrix_13_4 = 251'h67465ddf9e552984e871f6e16dced15270af54698a1c888db98f6edd65f7b16;
  assign mdsMatrix_13_5 = 252'h85a378fc9e4ae38fa9a4f1b9b905cfb55ca00a186b4bc23a574588c3484de0c;
  assign mdsMatrix_13_6 = 255'h4afa804dd6cea340257ecf00fddfd21cbc1d02d93af71c3399fc07588d6f992f;
  assign mdsMatrix_13_7 = 254'h2aeeebfff7d4d9848b68c4ad7cc1c5323bfa43a71c4826ee2376885af674f140;
  assign mdsMatrix_13_8 = 254'h2377f0d6770f3102de408567a0f778fc39ce39d7f37234b6ef39d51f788c25fa;
  assign mdsMatrix_14_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_14_1 = 255'h5ecb028cdc670317afdddc1f12a28500f5a24389d05291714eb18983da8dd71d;
  assign mdsMatrix_14_2 = 255'h52d02d37a509f50962fd3a8e7b51247e0c0f0fdf03ae3d85d3a1819029198ad4;
  assign mdsMatrix_14_3 = 255'h52416775390f7b191e74eb406a4f279870e90c81a7f199745b5fcb74798d2eb9;
  assign mdsMatrix_14_4 = 255'h58a36908f45a07562f2991f008000153178b95958e5cd98c8f32d36a96bde4cd;
  assign mdsMatrix_14_5 = 255'h66ee4759c262ccb642944ff6dfc69a2f2416a4f5f6b4cf5e94902ec6f45437fa;
  assign mdsMatrix_14_6 = 254'h3ee9ab84b88f634ecb3b9fe174ebfc49fc8a6a19bf89fa05805047871e79738a;
  assign mdsMatrix_14_7 = 255'h6c42f1a8d635bff4af805b13ed6a63d21ec8f5442731149f81dce6a85777dc80;
  assign mdsMatrix_14_8 = 254'h33bc52ab35b3484f5a5888ab69ff1fc591d66aa479a2b0eddfe17a1318597d28;
  assign mdsMatrix_15_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_15_1 = 255'h607442b4436c23ef6382f50350a1b9b73c8ceb026b497b0b16a1c3b6dc4a348b;
  assign mdsMatrix_15_2 = 255'h6d85b190325a58b23e8075c4a2dbc3514682a30dce554130bee5ac5efddf7c99;
  assign mdsMatrix_15_3 = 255'h54ea988660a5f94632f273d3613f79320698bcaa4b33b7f685812503e483bf7c;
  assign mdsMatrix_15_4 = 254'h3f2fe0cdc0e42f4455a4ceed936a8149dfa26feb7fafe90bb9cd80e3949c3cd1;
  assign mdsMatrix_15_5 = 254'h20dee0b6f58f125dd5cc3fc56ce4ced86ecbfa46ef289e2dd046d1176ba7861f;
  assign mdsMatrix_15_6 = 253'h112d5662d0ab0f9010af9086170cd8d2a223617fd2efcd91640a92bd10f5d723;
  assign mdsMatrix_15_7 = 255'h421304c4db679e65d0680f6d8edd2c7d26ca2a8f0190628501bf90fc5d0e83e7;
  assign mdsMatrix_15_8 = 255'h5599916626b57daa75a941ffd56daf9f8fa4f0d1f857fdb0572d2585c651d616;
  assign mdsMatrix_16_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_16_1 = 252'hf065f9fa6804a7fd7b67e04db743f1e160e20476e639589e9a479e2648e69e7;
  assign mdsMatrix_16_2 = 254'h35ffd2053ea9124d6e51544229df99419e3a319da6bbda1599674d50b6ad2f03;
  assign mdsMatrix_16_3 = 253'h1ee6e46f2308c37c308eaae837f329c72870a9cbc1376240255f0e688a3d4907;
  assign mdsMatrix_16_4 = 254'h200b65c292793ecbaf206b547e2e193410fa56a16e256bae10da68efa09a7972;
  assign mdsMatrix_16_5 = 255'h5dba4532b0f6a5157dbc463e0af623c87e0e9e1408f0a4cf9449cf3f1c928a80;
  assign mdsMatrix_16_6 = 255'h507305f8f4dc7077939bde862194fab4b2bc653cba27ab66cccc3687bd6c6974;
  assign mdsMatrix_16_7 = 253'h1f6418cc12cc98ef43e20a6c80ddb83002838097916ed487211214358c65c2e5;
  assign mdsMatrix_16_8 = 255'h47c162873b5f2ce5e08a72b0b2f6e1845ef96d32873e6a62f67795f9823a7392;
  assign mdsMatrix_17_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_17_1 = 255'h5f79fc6fcc6c72da9fdfbb4ec021fde9cd3d9cfade485bcf759cb120df9c40c1;
  assign mdsMatrix_17_2 = 254'h380f0e83ced9966a3050838241f8062d7d21e00644a8656390cc03b14d0d48a2;
  assign mdsMatrix_17_3 = 255'h5314e62c0dd570fee0a8feeb6f7957a2f58c05598975e764e32045bca554ccf2;
  assign mdsMatrix_17_4 = 255'h62f71dcdf62cd8d8b1dce4074a5f359cd02fdea59dada0eb8f2d163ba967ad9b;
  assign mdsMatrix_17_5 = 254'h2657705877124d1b8f2662b1c1c23fc90aec7bba5c6d3c555bf7ee25f3cf930b;
  assign mdsMatrix_17_6 = 255'h656578e2bf5f67d9be7a0bef42ab20a4dc39d9945e67c446e70338dc9c10a213;
  assign mdsMatrix_17_7 = 255'h5f17cca8b865806452ed678de95d12b485bbe7ac345f0f0ae1ff1dc12f69e459;
  assign mdsMatrix_17_8 = 255'h43db1c68bf98cf24b7327ab7b63fe2db4e39ef7474b8492191541f24be61e038;
  assign mdsMatrix_18_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_18_1 = 253'h11420dbff57918c190310f22c4b13d0b8ad32c6d3a9dd6c9e823856cf3b0f3fa;
  assign mdsMatrix_18_2 = 254'h24bbb3b973e324908c5b358d6f6cb444af6dc9ea2dd38d102fde1ab91b378d17;
  assign mdsMatrix_18_3 = 253'h1f6a7e0438513981912f825e770d2f9ffe23bbad27a7f5f09391ead2ccf949f9;
  assign mdsMatrix_18_4 = 255'h687e7a532039d2e03457baba079806a6a9576772278fee0ec102a2d3af89686c;
  assign mdsMatrix_18_5 = 255'h5df93d493d3d3445cac5dc5a5860cea4b54529c39b8f169b8e82620947068e4b;
  assign mdsMatrix_18_6 = 251'h6a6005930d767a24e10f96664abf1571280102d8a6ae086df36bf29a8a54300;
  assign mdsMatrix_18_7 = 254'h39db65769a6ec54fdef31e47d70f9c879e4389098d82662f21c82a5c084f7cdf;
  assign mdsMatrix_18_8 = 254'h3979a2b1e0bead3eac9d5a798228002c74099b112f8be05d4cd44b5c7b94deb0;
  assign mdsMatrix_19_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_19_1 = 255'h6bc0085a84feb6a415e09223a5b4c4db6824d5c63181bb4358b2110e25bf6ce3;
  assign mdsMatrix_19_2 = 252'hab6f524a440cb44912e535a539a0e9daf18d76eefc49ec35de064a6e1d0209d;
  assign mdsMatrix_19_3 = 254'h2e15cfc2728fd5424af8e818b8721fb46d0f4db54136304be9a1112eaa2bfe29;
  assign mdsMatrix_19_4 = 254'h3a7ad7762058d8f7a80748c31d8fdb6607bec6280c38847452a284dabfc48c9b;
  assign mdsMatrix_19_5 = 254'h210e705766465ae7ac115150bc6faa00160e1a8ea525316a6aa1484a001d7732;
  assign mdsMatrix_19_6 = 255'h662858a2ffe064a7b8470febe5ccdab4e7310590aca185ef349709cca2c4ea31;
  assign mdsMatrix_19_7 = 255'h7311c032d0e25c1d25f66d2e080d0ebabc19e8621f44cefe0fb1a4c67f174f93;
  assign mdsMatrix_19_8 = 255'h4cecbdde66556211d0b0e8365316cb2f3f7a97e4ccb4717e7143f18bb878f028;
  assign mdsMatrix_20_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_20_1 = 255'h4fb0b2020808703a54a00c09e05dca0dd6b812c1ffc7b35a633bf0e0d00ed45b;
  assign mdsMatrix_20_2 = 255'h603adfec029493481e40b358b3457517f228f93f6d9fa23924a46bb0b9c2fcb9;
  assign mdsMatrix_20_3 = 254'h330c1219b4616851bddec940a599a5d34b62bff7f32c528d050bd25f2d6db459;
  assign mdsMatrix_20_4 = 255'h4f94aba904a00fcabad13fcb146e0f7ec109e32478b4fde2d44257f25b2937db;
  assign mdsMatrix_20_5 = 255'h708a96d2d9d78ef5d0f7f29374a816772e9fe56d04ce951f97e7ce16abe3c979;
  assign mdsMatrix_20_6 = 252'hdc88a0341623a26417560a184d3a7af73e18adb046a1816121be9e73e0f5b55;
  assign mdsMatrix_20_7 = 253'h15fa3cd778461144122d2791e85ef565933f808f059b7aadcb08efbdaeb50155;
  assign mdsMatrix_20_8 = 252'hfdf0893083883820be10abd5c62d5acc15a18ba8bcd9ae39cf49309f49942c2;
  assign mdsMatrix_21_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_21_1 = 255'h41c2a7fab08c63f5fbd8d9af5786918fedb4b6a0ac2f77d990d809607b599dc5;
  assign mdsMatrix_21_2 = 253'h1f053429be53195620a18d4a471b3c96b1f3e2adbe4dcceec4e7cfc0b6cbb3e5;
  assign mdsMatrix_21_3 = 254'h2ba64f06f5f4ed1f2d2f676b58c385ebdb160fcc5d301a3a168d3dcfcaa7e776;
  assign mdsMatrix_21_4 = 253'h16b37cde38f3521d1dd4f5805ff17f89c32d75a3e1299e610547a44e2dbea388;
  assign mdsMatrix_21_5 = 254'h2148bdd4ce509a98050f444441ecf0a33ba16b79e1ec7c4a0846ca85a8d522ef;
  assign mdsMatrix_21_6 = 255'h4bd3f74d352ad6a027c4fe7d815adfed03511c773cc64613188acaee9ea88e73;
  assign mdsMatrix_21_7 = 255'h6aaad900d29f6888da0a34067f8921b2e69dee22e1b02de5419ccbadeb3600e0;
  assign mdsMatrix_21_8 = 254'h21ebebb0a1e023cb38c8a73824f7d66a2bca19495e92447609216e568477cab9;
  assign mdsMatrix_22_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_22_1 = 254'h3e8d82f4711d8529152523b9dc853c65fd5767909292a6cc6c706942f775c686;
  assign mdsMatrix_22_2 = 252'h8b70f948d28013df420023d24c65edc854d5aff5a4a55fac6ab4cbb63d3bbbb;
  assign mdsMatrix_22_3 = 255'h602cffcdaa7c19c389d02b75802e578d062d4f4e8c49d1049ef82cf71c9f37d7;
  assign mdsMatrix_22_4 = 253'h16322ea667f492b3c4081601b2ca193f66f1584e846255938204613736f4af87;
  assign mdsMatrix_22_5 = 255'h6098a66c309a79b556cb321188b38a5cb8bd7d2e7c2de719e39d88ed07a66957;
  assign mdsMatrix_22_6 = 253'h10b47769f40edc2cec2e86f169ef83b290c9d8b0066d364a55d1c6e47f0c456b;
  assign mdsMatrix_22_7 = 254'h3ebd8a8b412858ad6aad69c40e1f38c3722104ce09ab3ea0760f1fd8cecffec5;
  assign mdsMatrix_22_8 = 255'h51af1ca618e62926966c8ba0cd80e2b055b63d54b03a8d7964cc4cedf6888cf5;
  assign mdsMatrix_23_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_23_1 = 254'h26e1f22ed242fdb2f265aa2798f02bf15256150269abf84f02f2f92431654e98;
  assign mdsMatrix_23_2 = 255'h5262182f4a1d47e46583ba2bf795c65705eeb9f7e6eeed0ad4c1bbf53a37540c;
  assign mdsMatrix_23_3 = 254'h2ba0a5434e860abaad61a2ed2c7e6cff1638bca1e3e3e3ce0ea2f1ceed8b2c6e;
  assign mdsMatrix_23_4 = 255'h51c8735c399fec4d4f7f57c67fd2bfcc7bedffcd44e8da4365149567b6e21f28;
  assign mdsMatrix_23_5 = 254'h27a13845984312b35ef7bf6df2d4909fef1141a2a0df2763fa0278295beeefa4;
  assign mdsMatrix_23_6 = 255'h707f8ca2b7b1b275445b86aa19f186e6951a74120cb9fee2efb552f11d3456f9;
  assign mdsMatrix_23_7 = 255'h5b4038588f33959f26855db85a4d2b29f2cb1c918fa65fcd3cc33998488d8b68;
  assign mdsMatrix_23_8 = 253'h1c759bbbdc8e8dae10ab933c2d5c1329e59dc2cd10f35a2b39ac573800dd2748;
  assign mdsMatrix_24_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_24_1 = 252'hc36498749d72e13ae7dabee5d3d08e4b6314394d97e32403455fd96c50305d5;
  assign mdsMatrix_24_2 = 255'h503d44ab5cbd13ed7b0395d9435fd0c75b2cb39b309614a0f4ab0b57cf3b653b;
  assign mdsMatrix_24_3 = 254'h2fd2dc9128e73217a0597295df1a4c4e6c1e56f7c07f90999d903bbb2ece397f;
  assign mdsMatrix_24_4 = 254'h2d6e65538226389c75c627a31ac1a5da6ad98270dd7f919946232c491556b3d0;
  assign mdsMatrix_24_5 = 253'h187958987465bff067266f105f8033a5972149642714742382b7f34a48ad80ba;
  assign mdsMatrix_24_6 = 255'h41597a48349ae06aa9a9b5e47f2a900b93cd489fd6b00553e5d9e88251bd36ef;
  assign mdsMatrix_24_7 = 254'h30eba2b46a79a0009ef8eca18fc617686153199d93c8880a18f8fb1a34e6e6dc;
  assign mdsMatrix_24_8 = 253'h1094488e94b1296cd9a4e283e59b887b7213e2ddb6a8418387cec75ff5608b92;
  assign mdsMatrix_25_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_25_1 = 255'h5d437d93d385453f7ffa38d7cf74df4ea4be3b816268678d610d223e8f6a4c53;
  assign mdsMatrix_25_2 = 251'h62ce93688b36ae850c211c4cd4e969bfcc87c70e2c73ee5dd52ee721eda6f20;
  assign mdsMatrix_25_3 = 255'h676fd6393344a19a79367a01b1a5e00946777b68ef2f42010a78b611d1c34c54;
  assign mdsMatrix_25_4 = 251'h616767be41e6d5ed9f761427c89ac608a4659a3bcda07d14d1f6b3e086579c4;
  assign mdsMatrix_25_5 = 254'h31cf8c8ef4025ecc3e12140db4c4ca674c2f20575e2019927e8abc5abf82c87c;
  assign mdsMatrix_25_6 = 255'h676e7df1b170c51e088415f2ab2e66b9432d2e8c846484f584f0c0a22aeb6b4c;
  assign mdsMatrix_25_7 = 255'h55cfaa984fe0347abf9101cc326b39bcf14cbc0b51be80c3b16a8844adc5f383;
  assign mdsMatrix_25_8 = 254'h3c4615a20d1901686188c8ca6d7d7db6cd42235c7c96d841a7df16b58843c8ba;
  assign mdsMatrix_26_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_26_1 = 254'h241f111d5623012b2ae957734a27c08c2636d4e4b4737503fb3225d79025c3c2;
  assign mdsMatrix_26_2 = 253'h1c7d88122970541aa6a4ae241456044e83d2c08ad93718eb975659e25f221bdf;
  assign mdsMatrix_26_3 = 251'h597c59911d9d0caacc5b6366d8e23a1ddb003cfc0e35df3b16c9fc70e6f395a;
  assign mdsMatrix_26_4 = 255'h5c92d0fbd709e67f27437025f7d37e93f32c0cada03d402085ec6624568ad03d;
  assign mdsMatrix_26_5 = 255'h5400907800c95b93fffb031b46d7701da26d3a21796d3321978cf2b891e98804;
  assign mdsMatrix_26_6 = 254'h3f6567c993eeb9e8d7ef7e62a7011fa2a5f1cfe86203ecf40b7c8ba2e05b0646;
  assign mdsMatrix_26_7 = 254'h325d69c0b6c794eb87f46af0e3c61a25ae1516fecb20571aaadcb826f36e54ee;
  assign mdsMatrix_26_8 = 255'h5e94711739fbbb2c9a6c53ffdd7abe082d1f5bfefeeedadda9380a3e02930b16;
  assign mdsMatrix_27_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_27_1 = 254'h2cdaf67a16f52c87bb003801aa4119eab0940b5c8353ed813e0d740c0f65d9aa;
  assign mdsMatrix_27_2 = 255'h5e6dddf14cc7f4bf7d70255da91d11e721cbe217f8f20669956e5d215a91d75c;
  assign mdsMatrix_27_3 = 255'h6450ed3bc60c67c9a99e1153ce129fd6400021d6c4a186c2d708aa7db23279ac;
  assign mdsMatrix_27_4 = 255'h4cd61bcd82d3ce386423d96cf6abf3c75b3d5191528a100879479081699a44e8;
  assign mdsMatrix_27_5 = 255'h6f11819e593186b739d6cb00827d00e8af2f11abcb0417ba26e0d0ed1eaeea72;
  assign mdsMatrix_27_6 = 255'h66ba04c4fdc294820ce779ad8aa6d47052a64586b0cd431922c864a01cb2b64a;
  assign mdsMatrix_27_7 = 252'hb9f59e78cf286504dcb5d947380a9dae9e9c41463b95349bdb70c7fe06b3dc0;
  assign mdsMatrix_27_8 = 250'h242d9056a66e36c51b57f8c2d6c063e83b04ea8f74b5f64d835bb02375a0e58;
  assign mdsMatrix_28_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_28_1 = 255'h7218ba28122b82f709ff273f2887dc81a54be5a500da09b6cac81531b4019e0b;
  assign mdsMatrix_28_2 = 253'h167db00df9f6c2a685582250d8bb40756a0293dfa694d6dfa4f9ea74733f0b59;
  assign mdsMatrix_28_3 = 252'hf8094dde36d9d9121b8d85514ef62e110de285a9cb6e739bceeea6c2736219c;
  assign mdsMatrix_28_4 = 255'h5e63a054ee4eeff069ff151b837e1c84c0293dae5892adc730c9622f379cfc9a;
  assign mdsMatrix_28_5 = 255'h73b30ad2354b23601e1f787bee546505cbea80e130b5f975acfbb73283b2c678;
  assign mdsMatrix_28_6 = 255'h7160a2238a75383bd85e77090d3a2df40cd8aa2a9272c5db919d35bbee11d622;
  assign mdsMatrix_28_7 = 254'h2ecf6147404cefa4b42b1371179c5d00eeae5801816279d1efd8a25a0add7a33;
  assign mdsMatrix_28_8 = 255'h70706ca64731e35bc93cab846f01f0dd6fddebe6af1cf86aca7d56e858293f7c;
  assign mdsMatrix_29_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_29_1 = 255'h65ba89174411b426ab118718794f51d3c8c961beb803fbd52094d0c218e66ffa;
  assign mdsMatrix_29_2 = 254'h2e2e33043873b29e8b538603ae3a3df2929cb741f5e736cb30cad345c385fe85;
  assign mdsMatrix_29_3 = 255'h48cfe06dad8096f82ea8c68c692de604308d58dba83d55d5c8bb8f40c704d87a;
  assign mdsMatrix_29_4 = 255'h6d752b00b38df17771fc6aaad8326f3f7eb28057f8f45aa2b17f92bbe849d8ae;
  assign mdsMatrix_29_5 = 254'h289cfce097541802f8b833d3b5a811a2e4e7dad4bc673d4206d0bc54380e71f4;
  assign mdsMatrix_29_6 = 254'h2bb81ad56732ee46c126f6b8845c4bfe6ec5e2a645c5ad4d3a268c36c91723b1;
  assign mdsMatrix_29_7 = 255'h5e06bbcf8cad21d759d269c11a07527f9fd29a292c14ef3683ef52c446d2b6d3;
  assign mdsMatrix_29_8 = 254'h39c2e3437a0b18cf7dc941b61b9ad7c4d8d71bec2d5c0de92f2ec77709e34f6a;
  assign mdsMatrix_30_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_30_1 = 254'h39d3ed4d387748108fefdd5ae3b88e8cad4519b14be1c0311bba1714cc5969e7;
  assign mdsMatrix_30_2 = 254'h26bf740cd9f871c59860d9f5cb1249c0da9485e487d98b68fa982e4722cd1115;
  assign mdsMatrix_30_3 = 253'h1df57e15bd844384ec525311d5c9685d24f1ef3704073f26d05c5c90551f0c05;
  assign mdsMatrix_30_4 = 255'h63e0eed973dc8a38051576f493ed44da17598c10c540a5684fbbdfd7c4e5efe7;
  assign mdsMatrix_30_5 = 255'h6ee4ef50a40382b4f67a9a976156b5364555b4d9db15ab66e7677e9975af574c;
  assign mdsMatrix_30_6 = 255'h5b919d85727f9eb38f08d5033d9a41d6b2ea40fcc06587d47960b3907d826963;
  assign mdsMatrix_30_7 = 254'h39d80eff7b82a94719583d4dd1e6ad84c9e127573c854558245527b2b2475de7;
  assign mdsMatrix_30_8 = 253'h1b8b0a37a095ffc8d3a4722d109f5ec91b9a5966832a44e90dc2638f5781f411;
  assign mdsMatrix_31_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_31_1 = 253'h193734b9a79c9cc8bfa6bde8d6f850c515b1420387ed16fb524c79e223dcdc0c;
  assign mdsMatrix_31_2 = 254'h26cb29a9d1a69179436b206abd86022afb50a7426748b19f96030da50d5e8c68;
  assign mdsMatrix_31_3 = 253'h126c6f710e17f29f583a3d8adbee5cef16e6857662b0048c8b9940b6501f97eb;
  assign mdsMatrix_31_4 = 255'h63bf1d5d20414642437ca50ec8262eddd07af7f2605051821b5c58a2f1d2fc09;
  assign mdsMatrix_31_5 = 254'h26d0d3b9550700196c476f70738f5b52df0409a66dd45cf85b88f10184adeb6b;
  assign mdsMatrix_31_6 = 255'h40a4d203414f89d8f8c543e1eb5bb67ca5bdb4a3aa5d9a6d2ee87eb1f4b19adb;
  assign mdsMatrix_31_7 = 255'h5bdb26c8170cd9386dd1cce66813aa0b1edc81fde438a8be28bf571c3f594673;
  assign mdsMatrix_31_8 = 254'h241f26b90a0e97697f950d8a937d941c72b1828eab7ded74a56547f71731bfcc;
  assign mdsMatrix_32_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_32_1 = 254'h21bf2e10c108b29af050bfd6731dbcb52dc28faf1acda962ec1c64caa3d2b358;
  assign mdsMatrix_32_2 = 255'h6797722155f7717f23512f0f65452c1ae1610f031bd7c36d8b10ddc1a74194e2;
  assign mdsMatrix_32_3 = 255'h60b1f1bcdb3c9722329992768357b053260bf46546177f2c66ff3c1fcd648281;
  assign mdsMatrix_32_4 = 253'h18fb82cc867d267ce18fa986f17a1438c281223f63f782c921db65008d67c814;
  assign mdsMatrix_32_5 = 254'h202eac98ffc67347db7f8ee47263380aca7425a40a35bf80002f4d4ce250a1fa;
  assign mdsMatrix_32_6 = 252'hcffbe8211c00e557487fc2769dd2e27144544130fed7ec3fb7d66a3f9c6b29f;
  assign mdsMatrix_32_7 = 255'h5720c88c7453a1a5acbcf15c207f6fbf778a1318b4e598af3f6102cef66700cf;
  assign mdsMatrix_32_8 = 252'h8b17bbee1b6b6d676a366248f23135b6d42e23a5f9e97814271c39949c16bec;
  assign mdsMatrix_33_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_33_1 = 253'h12218dd0eb67d9efa4f4d7ee99fe6a88b665652d96a91c9878810af4f6830217;
  assign mdsMatrix_33_2 = 255'h58fa1f3d7b0cc59a86e66e425634b517b83633db3de41bac760c0d488167067c;
  assign mdsMatrix_33_3 = 254'h202e71776d871f9a0188d5da15e3ac80aa69442974ec92caf7e7e3e3c239d543;
  assign mdsMatrix_33_4 = 255'h4e1a0ed620e2f5ccc56e9cfb52d387c16c17e6e8e68b9f82ee13e2b47c41dbac;
  assign mdsMatrix_33_5 = 254'h343dba558e2619479d9135e0fc80b699ac4e958f68046110908065c0036c7d3a;
  assign mdsMatrix_33_6 = 253'h1d6e974ab405e28d0f2a79b342059be71d610c68aa5e75014f853d2c6e038a2a;
  assign mdsMatrix_33_7 = 252'hd675ea8e29563628577885cb6b7e419dc1e657d3e9123069c10715f30495142;
  assign mdsMatrix_33_8 = 255'h5e165278c8f1df014ba1bf4fac4283984e44b5e17c38a9ca08082bd354c35f24;
  assign mdsMatrix_34_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_34_1 = 255'h58d67290655e60018e8c0a805f1eedf428d6cb468cd860733985c2f9f1d02ad9;
  assign mdsMatrix_34_2 = 253'h1d9eafc057bb4953e80a330de513e079284590b0eb75ea3d7735c0e3e3c6ba63;
  assign mdsMatrix_34_3 = 251'h57f11c500f0ebde02b035085e56acd8073bd2ec3f3ee274bf1f43cb5e8bcbc8;
  assign mdsMatrix_34_4 = 255'h5cb19435b0459712f51f742b317d843db344359e011cdbfcc8bbc23529848428;
  assign mdsMatrix_34_5 = 255'h591ce4f71c0b194d0e29bd16ea381a4e39b87826730e618278588964fdcf2e16;
  assign mdsMatrix_34_6 = 255'h4e895a57c8374eb11180dc37e64900534a009b16a9a7f5a8d752e3bd7e29f4d3;
  assign mdsMatrix_34_7 = 255'h6f408d731e364ffb9682453a64ed658de203f2f868c0055dfae7b8b84751e665;
  assign mdsMatrix_34_8 = 253'h1df46fa8203e5db5bebeed90b8a18e1547ad1f0ffaae0d082be53eb01dcf17de;
  assign mdsMatrix_35_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_35_1 = 255'h4ea5b033fb4eca2d5c9c02f9820423c588e22ed483f3624e7d5e9c3e0f9ad287;
  assign mdsMatrix_35_2 = 255'h68b7dac95da1d73e63953d9dbf6ff36fbcc5b847e980369acc5dadc8e4487c48;
  assign mdsMatrix_35_3 = 255'h4df8871e093b3c481c889d62f84316f527189d9895842a6fc193bec17f5fdf78;
  assign mdsMatrix_35_4 = 255'h7305143148907d27a2debdb3fb11564c2acf384a1d86a9d02d74a0a194836e17;
  assign mdsMatrix_35_5 = 253'h1f3bdc57a6b4a5e8e18183f88fe3a1516ec9650011c448d64fba5f68cdf81e20;
  assign mdsMatrix_35_6 = 255'h63d0fbd793af05270a6e4fe30bdb45cc5594c0113a37e8227d7486236aea6252;
  assign mdsMatrix_35_7 = 255'h46e1ab3b22109a5cc0618ed06b3c25da716e48b72969a2bc09a78c58a8fe4326;
  assign mdsMatrix_35_8 = 253'h1cd4272b216ad0717150036bbe88dea602a0d5101c4bfa16ac6ffe1e2458319a;
  assign mdsMatrix_36_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_36_1 = 253'h139374d30cb1fed988757f7289f1257da4be5fd9afa854c28ad8b81c7afaea01;
  assign mdsMatrix_36_2 = 255'h739d79df930443e324bbd19e749af4274cd2f01d97c5efb94fefea46419e967a;
  assign mdsMatrix_36_3 = 255'h4e2c4d00b708246ac9e5fe36a3262655ad7b2e66f50dbe10eda16685b26c24df;
  assign mdsMatrix_36_4 = 255'h61752d43aab45ac4fdc5e681fec7e47c3bea42a46dd4d24c5d09f99e4dfebecb;
  assign mdsMatrix_36_5 = 255'h403967e0c5521951d61ff93e424d25366e4551e9872ff479f9c81f945e5b0bbf;
  assign mdsMatrix_36_6 = 251'h66fb6d21040e9c609f53be750ff8cccac2d18df1f2d9142a447c71412862339;
  assign mdsMatrix_36_7 = 254'h2ce5fd6c958e6daf84b4e1b0237f7363615f52e3d2f5bf067c922310835ac7c6;
  assign mdsMatrix_36_8 = 254'h322eabfecd954e0c2e85eaad799f63b67ff50cd45ec6c584025b576115d56e19;
  assign mdsMatrix_37_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_37_1 = 255'h64d87f5d21e519cb32d58170d695aa264bc556d42eb6cd679e6eef069909508f;
  assign mdsMatrix_37_2 = 255'h6554cb810659721675d7cbf63abd1842805f5b4e2842d0f0875e7dd617dadaa5;
  assign mdsMatrix_37_3 = 255'h5da01a44c7f9ee81462bc536f5ff58d32f9be08c110d13beb1cf0a1ab9570090;
  assign mdsMatrix_37_4 = 255'h575c937ea16964132885e4070298ca844084a70906550b0ebee941568050a521;
  assign mdsMatrix_37_5 = 254'h32941de274ad1f8acbec8f5d3429835c8099cf8e5221cc2d681fa4d92148c8d0;
  assign mdsMatrix_37_6 = 255'h53cf4eeca3439c5ce98210ffc0a8e04a8ee4245698789502688e361086cc9dbf;
  assign mdsMatrix_37_7 = 254'h2e1444c94a7f93c9c11eb6ff81753801537b45ed6cf45f78e3ca9e22ad7db8dc;
  assign mdsMatrix_37_8 = 255'h4bd7dc106f1769e0ec8f3dcfe6b484f650c880b2e289689e2ee4ffed4443085f;
  assign mdsMatrix_38_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_38_1 = 255'h50702599d49b874194c7ee2a6238d600d358a719a4bb3023f7995e767e908b1b;
  assign mdsMatrix_38_2 = 255'h5baec648b50d64128296c517090a6464ad25cef403807a35d2a50b61287f5068;
  assign mdsMatrix_38_3 = 255'h4121098a3156f76f0d79fff20f2c0fa832658b4464b6a6480f559f4d86130e6f;
  assign mdsMatrix_38_4 = 255'h499225a97c302624437687c2e54894856c124548900238696605af98bbeea844;
  assign mdsMatrix_38_5 = 250'h2c20ac95195e46b62f01a24e074f0a1722c98f6306291deb07f0978d6d1a33e;
  assign mdsMatrix_38_6 = 254'h2ffb1ffaa88f7761a21a1a750ee6216abf79e5e39173abbcef9a2fa7df1f0a6b;
  assign mdsMatrix_38_7 = 255'h65bcb355c0a39844856f8f3f597eb2def084bc9766275624ced5c0da92fc6ecd;
  assign mdsMatrix_38_8 = 255'h6efc7385b772973fdfc59f9584b6fb16bfb11f7c54b5084c2776c51ec318f425;
  assign mdsMatrix_39_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_39_1 = 253'h17189106174ef9fdfc54aace80e20e55cfe3873e1873dc9b4a9a20b3980ff157;
  assign mdsMatrix_39_2 = 255'h4c05066e28ade8ca7a36c4ccf551cbaf9cd1b2320597a8ed422987c2b0d208f9;
  assign mdsMatrix_39_3 = 250'h3dbca2407fde8a73b222e973b507b7250e6106a2dc1674a4fd600952e5192c2;
  assign mdsMatrix_39_4 = 255'h7036e553b547a5fc0d59a3b1c83c77b6de06a04c5ab52f381601d8994bfcb739;
  assign mdsMatrix_39_5 = 255'h6d2981726f619aaa6e430da581f43151ac54f7843bbdf73a028c9ab53bad5ffe;
  assign mdsMatrix_39_6 = 254'h3745d0123f9153f0bc0655f3fd4f48a9fa53cf0d714dbb3b1d8361cae6d36975;
  assign mdsMatrix_39_7 = 255'h584cb1e18736e0d56f85f332ca670ef4b6fe469b2a99448cf2ec61f4dd83b74a;
  assign mdsMatrix_39_8 = 255'h51d1d990afdad506fddb2a97acc3e80161cb8bb92b59c646e2a40192a4e3410a;
  assign mdsMatrix_40_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_40_1 = 254'h38a8b1a17861641ee9bf23557b034e48af33f5f9de1db1e5f5b1e26209d48105;
  assign mdsMatrix_40_2 = 255'h4878eb4e59b2ed4a29ce48282d942fe7c08e8738707f24bb3eda9d76b48ae46e;
  assign mdsMatrix_40_3 = 254'h33969085822da986a28b313a86942a141cea96d6f9589f7274a853316231f714;
  assign mdsMatrix_40_4 = 254'h3c126418c6fedbc3c84b3c5462b5b1258bdd80c2d27e8c4e6a9649f64aa72997;
  assign mdsMatrix_40_5 = 255'h665f04a97d1a824c24eb331640c2b9bf7e3f3b75c3b96a1ca5dc7b7c2f4af132;
  assign mdsMatrix_40_6 = 255'h606b643015bd32bc0becfc342b232a20184775dda1d06c226b73960a389b9966;
  assign mdsMatrix_40_7 = 255'h628bc43bf4b560df7732ebc589a8bb2605de704183573e454bc0b17310c9a4f6;
  assign mdsMatrix_40_8 = 255'h4520ae8bbe3317e7f4177dd14595905ebfb0f35ce35490f3fdd4561c7fcb3f8b;
  assign mdsMatrix_41_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_41_1 = 252'h8aa20c54b37a2d09ad1933c912dae0b84409080571134b5e7394ed7c8381aa3;
  assign mdsMatrix_41_2 = 254'h296f2352d94651cf5d423a2f8f4bd62cfa161fdec7a176ff21b4ea3e33a32c7e;
  assign mdsMatrix_41_3 = 255'h67d1012ef53e49574ed53a0bd1359da157860eec7caea6b6a96ca00472f45786;
  assign mdsMatrix_41_4 = 254'h2f9020db69500aba11dbc5ffa7749a9471967fc3c92acf54590212a3a89231df;
  assign mdsMatrix_41_5 = 255'h4dc0eb99b8937f566f1b8fc379bd6460c72ea570a5aa14c716fa030f10b15143;
  assign mdsMatrix_41_6 = 253'h1da2f8de49de9b9ea1d0d93b23a38f7b6f2ab59cce6116316703ebd89262fa9b;
  assign mdsMatrix_41_7 = 251'h68504c2b606abc5245ca724892a29dcad9ab00352e84945b61c36e0b1143d02;
  assign mdsMatrix_41_8 = 254'h37422ba9509cc61aeecf4fd751f37f8e6219b913a30e08d650a083c7171a9177;
  assign mdsMatrix_42_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_42_1 = 253'h1bdabe021eb58d41efd3a54eac47eec3f4c52a874543abf857704dfab339489e;
  assign mdsMatrix_42_2 = 255'h55bff0893d72ee0f7f4fcdfb79e7342328b153979b2a7f5cc9f8ae213d8d6e78;
  assign mdsMatrix_42_3 = 255'h49b3701dd5dde22a7bbbc90127099cc5fe52af9bcb7d547748c3010fdecaf6e9;
  assign mdsMatrix_42_4 = 255'h6ddfe17d9c3b4f30816e5662a041fb363c9e141a012d06f97f080b31f0358941;
  assign mdsMatrix_42_5 = 253'h15efc155ca424cc5ea76ccfe4a4e91956ca7158918b2056767c88f914db768b1;
  assign mdsMatrix_42_6 = 254'h27628a2900a0dfef10109ad08eb7d9b11ab279b2e68057063a16dabaa4bcdfcb;
  assign mdsMatrix_42_7 = 254'h37da675b6077fbd1fac68de30e6c07344af1345d983973942653ad10b2cec6e5;
  assign mdsMatrix_42_8 = 255'h5655761df168b518cf9c3d60edf2111fc19a072d145078fc675db3e8ce6a18b0;
  assign mdsMatrix_43_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_43_1 = 255'h5282f727dd63ebd6acb66581ad767974735c6932eea147c9d236f91228609de1;
  assign mdsMatrix_43_2 = 252'hd06c6e88f1882923ae664f419052447bf3f9454040431412bd12806f62d08d9;
  assign mdsMatrix_43_3 = 254'h31cb729bd1fcb0d3fdd5797a597ffa9f60abe6e8a7a689f3e1c3a9d7c6e68a1e;
  assign mdsMatrix_43_4 = 254'h2a98d712b49e701c56f5eeea650f91d7da8c0500eeab5b8557a25cc9430a9e54;
  assign mdsMatrix_43_5 = 253'h1039c8798a3ce13e576094379c82b0a847301c7e110d212037ade8c7843ddbe1;
  assign mdsMatrix_43_6 = 254'h32710ddfc5df75ed86bb86c7394c049e328ff5c9ada2eda178d5ace13a120ea4;
  assign mdsMatrix_43_7 = 254'h3b83fe1083e763e2952b2dcd6e28981f912c4aa2f04e1916368576d8161ad31d;
  assign mdsMatrix_43_8 = 252'ha3f0def6f657f6c7a8566a46dab3c0ac423c9d27a3aec5a5113d8407df0c2a7;
  assign mdsMatrix_44_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_44_1 = 252'h9a3654e2445e13f69334c4aeb6a3367ab0c15a863ff1d44389361cbd2389b29;
  assign mdsMatrix_44_2 = 254'h31948c89edd875febada7ae677f258b7a3320deaa1c4c5ff826dfb5c4e076f8c;
  assign mdsMatrix_44_3 = 253'h1d2deaa87ecfdda948bb39b2f92288bf9217a00b45e86d077f914f0e5d7197f5;
  assign mdsMatrix_44_4 = 255'h5efc3e2e0a522c31e9d9a130200542bbd68ce85e27884dfe6652eb33eb4d4895;
  assign mdsMatrix_44_5 = 254'h36890f2d3c8d0b730441bc98fde6bb7ef51021d0026a0f72afb00cca980848b6;
  assign mdsMatrix_44_6 = 255'h44c31be0a29afbd898123d29f6b85595b58845e17ef6b46634055badadf38124;
  assign mdsMatrix_44_7 = 255'h5ee7bf93d16320afa59598ad88367561e5b8bafa8f36767754ac85a5b71d3dd4;
  assign mdsMatrix_44_8 = 255'h67fb87fadf6b05b2301e91b5e202216bffc0f6ec345f808a00b054a7afb9f13c;
  assign mdsMatrix_45_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_45_1 = 255'h6f2b02608b7a1bbf172bd9d1f361da30fd1082a1e4ef294b7b5a000846c17dca;
  assign mdsMatrix_45_2 = 255'h47bdff4a8e90ee4ab6d3f11a24d3537ebb3e6c6eb767cc1b27854a1411d75fcd;
  assign mdsMatrix_45_3 = 254'h2dbf48ffdebc507ec4e5ed2c1607361960e679e0e27d5e698b497492f1131023;
  assign mdsMatrix_45_4 = 250'h2b2b2de87aa84d75368aa7ee00592c33fb4cd5a61845288f243f0bc83496790;
  assign mdsMatrix_45_5 = 251'h63b28739c793034a25e4213a58d5dd9814ee45ea40bd8e04f12547375d9ef43;
  assign mdsMatrix_45_6 = 253'h13c231fccedc7613f1da58dd72ae9586d072b411018e85973387136669f9e007;
  assign mdsMatrix_45_7 = 255'h6b83a40950e2e28e38bd82a88c8edf5276b617324d25ed6bbd70891a9e47ff87;
  assign mdsMatrix_45_8 = 255'h4e781e36d2b5a7d2f99096e937548ff938dbf527e505eb106a2d605cf5f225eb;
  assign mdsMatrix_46_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_46_1 = 254'h2c8fc5605cad910a08c995150d968827507ef1c2e2648ed6d17183896a2e5d59;
  assign mdsMatrix_46_2 = 252'h829ce63b5e4a6f823b9f0d7a0752f440166cad794afc6806882f15da2e6bd89;
  assign mdsMatrix_46_3 = 255'h4e39fab2fc0c3d9e246eca0c31dac5372ace1aa4444da7aa52b6b369aa271039;
  assign mdsMatrix_46_4 = 254'h3f7e8f19262d300dd13325f1a5ba78a04a873d4f4ac305e1b477390a232f944b;
  assign mdsMatrix_46_5 = 255'h5edf408fdf9534d3f5b31b7624f49839fa38724eafc92d945b75ea819de703a7;
  assign mdsMatrix_46_6 = 255'h72be6039f27acd31251ccf43e096efdfadf5ae3e4d1240040f913a52a9086383;
  assign mdsMatrix_46_7 = 255'h52dbe7bc46453ab761711c3a15664c3fce8666c3aa68d8133c90e2a8f5ec1ee7;
  assign mdsMatrix_46_8 = 255'h4848f5908290fbad9c2742c0179480ae7d13d674bff3975fcd2ef11ffd67bf2a;
  assign mdsMatrix_47_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_47_1 = 254'h3fd7a2cfc1842674b631df432d4bc4fcc03bfa130287ebdbd29a4a2a65a9bf46;
  assign mdsMatrix_47_2 = 252'h9f606e31dd715828a87d780089134d403c984b3054f026f8e6a589b7cf1beef;
  assign mdsMatrix_47_3 = 254'h2a9f93db8e3d05ebe47470f393c7e52454153636ffc1d9038d3f44f40b97459e;
  assign mdsMatrix_47_4 = 253'h14e1e9869fa5dcfa1d5bad76ff7cba746560d9cb6e782df06b80619b90172464;
  assign mdsMatrix_47_5 = 254'h225933f77f7b02303c0b098f7d21e2dcee85a24c5d1796fb4eeebffb08e298f2;
  assign mdsMatrix_47_6 = 255'h6e83fd6f8edd10e46f70a3e015459c7a414c49e3549c9bd383493a554e21d382;
  assign mdsMatrix_47_7 = 251'h61024f06377a17b1179af6198ebb1db3cd68e6d37a00f016803346b468d4e19;
  assign mdsMatrix_47_8 = 254'h2649cb5a8f029a2a6eafcc0079f2a5f0469ee17942eafdedefe43baf3ae15221;
  assign mdsMatrix_48_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_48_1 = 255'h6a4c66c4d54672a4d9777b25c576b4e6fe6f42783e9c6c77f218003ea6a7a2c0;
  assign mdsMatrix_48_2 = 255'h6573b39fab82f6d0f7a29db39628c244a84252de2faec0720d03ec857628d04d;
  assign mdsMatrix_48_3 = 255'h568ff17afb0d8be89b61ba61018a42686af75b02173c3c5249ac8dfc4a681240;
  assign mdsMatrix_48_4 = 254'h2875020bf45adfc0bef21ede53cf2b722f91c81707eadfa148354fa58fdc9c25;
  assign mdsMatrix_48_5 = 255'h62359212465bf41b87b327f2ae9af7408b133c0e39c5ab7f995743f15088ccdd;
  assign mdsMatrix_48_6 = 251'h74093728905ac64c4b2bdb9d95cbb203f08600cd4ca226c38571b0de8e1fc7b;
  assign mdsMatrix_48_7 = 254'h2b2469b512863d0383c88d5caa6453daa78aeccddfe4aeaeb5ac3d77e9744bc0;
  assign mdsMatrix_48_8 = 255'h5f189500e965baf7d5cc0965821979b620b8eadbf55d4cfcbb8a57e8f7b9d38b;
  assign mdsMatrix_49_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_49_1 = 253'h1195e866894e57ad209cccc1c76c5020319b625d6e6ffda5188ec4a3f2faa7c7;
  assign mdsMatrix_49_2 = 253'h1b0a149da9d17d1b273e88f31da389a1ff14ab4689bf424f93862828fc0a42ec;
  assign mdsMatrix_49_3 = 255'h64f42e5eb80ca356f196560f5962aa813b447245b8bb5cc03b6b4e5620c2bee1;
  assign mdsMatrix_49_4 = 255'h5b6f3a5bfa22d162936dd29b2b514c29554b9ffbc29073874a38f0929f5972c8;
  assign mdsMatrix_49_5 = 252'h98112aa4835c61e877a535979530f493d48b074ab53a5cfa8c3b4611437522b;
  assign mdsMatrix_49_6 = 254'h351ed90d2091798dd9ed5e3ddaab4d53303a2a6f3417823d876017a1f07377c6;
  assign mdsMatrix_49_7 = 255'h41d0c22203289e0a6f908fba41af5040d9d0bd06188980f08509c785ca3b9702;
  assign mdsMatrix_49_8 = 255'h4d68b474aa9966204b5e320ea8b889d39afe2e472c8a2569e1ffc7804889e771;
  assign mdsMatrix_50_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_50_1 = 254'h3eff3ff20facb905eb909f2131d61993696c51533410e163c9067a9fc90c7021;
  assign mdsMatrix_50_2 = 253'h17356a4ffb232c311853018050180243005da6500e3f1e3a8887011818ce785c;
  assign mdsMatrix_50_3 = 255'h66cc84d147a7455fddf84b2f110248ef4b3417620316f597ffb4666714749d3f;
  assign mdsMatrix_50_4 = 255'h43c1d3c719cb930776553515576ec6d87b43954b5e75fec69bd01537968e85e3;
  assign mdsMatrix_50_5 = 254'h302b59d1e1ce036e1642fa0c1c8fa96e0372774f71a51fbedf2ccae78b29ef6f;
  assign mdsMatrix_50_6 = 254'h244103e59fa87bbae7220a67cdda358f295f4d7f8341db2c8d3a13e2380fbe5f;
  assign mdsMatrix_50_7 = 252'h870523c2258bac6bf2b94e0a84ba8d62f35005c9eb49cc10c044c2ce1655167;
  assign mdsMatrix_50_8 = 252'hd7d53550f3f5c8dc1e6d4cc57bf8f3aa7aed5b9878719824e3de50fe91f2f6f;
  assign mdsMatrix_51_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_51_1 = 252'hf8091bd1d2f23f27764be07071888e6d75933c5f39b8aea48a5dff5928ba205;
  assign mdsMatrix_51_2 = 252'ha811bd00c67b4470f17fd2f109ff2386656d874b1dda15a6e8df7359084a2fd;
  assign mdsMatrix_51_3 = 251'h4b71a1eacda727c3ea4b63903145d7db33e3e0c7d577c490e09a26f7e8ec82e;
  assign mdsMatrix_51_4 = 254'h2c50dead0d8377ad7bab332d1b9e461951997119eec2acb618ae035cc5d60c9c;
  assign mdsMatrix_51_5 = 255'h6423cfc4a1ba8db73a46dc2d930f027a00b881cd5db0d60ea8eac6c349ec7b18;
  assign mdsMatrix_51_6 = 255'h49cd3945a9a3b77faf57584de3d115fe2719967d95ae3e7cea24463bde6114ce;
  assign mdsMatrix_51_7 = 253'h1649388684cfb6f4ea72baffcdd518e702f9db557291ab40b459c58d72413c3a;
  assign mdsMatrix_51_8 = 253'h1a3e37c5dbdbaa4a4bf25e28bbff4402cad141acef20320e6fb23482a73a81c4;
  assign mdsMatrix_52_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_52_1 = 254'h2ef34fd5329fb9b0ba7252443f1a0cd968ca74bab87ffe3c3637b1fd01cd0514;
  assign mdsMatrix_52_2 = 254'h3b87302e66e65d85688d134ecd2327712d2c9966a6bd6e20a9b996fcd448814c;
  assign mdsMatrix_52_3 = 255'h6124edba1994795198398261521dd20c08c001748fcbdef1e748d8f588dc6635;
  assign mdsMatrix_52_4 = 254'h3121e1808038653ac472b7b15e17a00fee19031532e6aa5afd079690f4f3bbcb;
  assign mdsMatrix_52_5 = 254'h2850f74d9384ec81df2897a764f6e38fd8e68a283a45d6875877b5cf4d052d09;
  assign mdsMatrix_52_6 = 252'hc7379c23812a8c37d71c77dbf6d1c9a8f49ab24dbba8f288b0fa1426053ac0d;
  assign mdsMatrix_52_7 = 255'h643d4fa266da84460a6613850e0063a5e8918b9a557428f436b2c92974514fa1;
  assign mdsMatrix_52_8 = 254'h2ee4741bb9daa2a7408dcd94f6e4b9fb59c227d6be2a470e5a80678ab03bb740;
  assign mdsMatrix_53_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_53_1 = 252'hc79a6a82e250192451921e8d65dd2a716645ce90612f43ed2f3f8f1efdc573e;
  assign mdsMatrix_53_2 = 255'h5c8c43e53277d21a6d5218e7f887471d68de5831f4233696311e711b37d42201;
  assign mdsMatrix_53_3 = 254'h37fb21180d810c8cf5eea2541951b9b49f5ee87490d7d6b74c3370b36fc49432;
  assign mdsMatrix_53_4 = 254'h30d72bd2442469c574a206611f4bafbf39a3b6306872cda1824da8303a64dac9;
  assign mdsMatrix_53_5 = 252'h877bf0877fa65fc4993536dd81030295123703182d7b7ddd6169aecd4934bf0;
  assign mdsMatrix_53_6 = 255'h47ad67bf95ebce34684c12765a386ced5335bd014f2f6dd201ad79f3fe55c21d;
  assign mdsMatrix_53_7 = 255'h6894319cdaf73881fad646fa45f123c5bb1b1853ce2cf915312df4823c8480a2;
  assign mdsMatrix_53_8 = 253'h1c75c65abebfc6923da0c295d0e9a01f6a300eeff78c28e26e3248210fc7876e;
  assign mdsMatrix_54_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_54_1 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_54_2 = 255'h44ae2b4dd47a8c0b601e049b50781fa47b173c9d6c28e982f959c4276f440b87;
  assign mdsMatrix_54_3 = 254'h3e392f76040ddd0f9b1a70686f9af4355b5d7385b9e2341e50e682c4d8664093;
  assign mdsMatrix_54_4 = 255'h4e55444bbe4e5727e8bccb3cadacaf2dbf8f78afff607bbef61c790cd0cb985d;
  assign mdsMatrix_54_5 = 255'h46510732b4340c068bf03af067a7e48373a7df79ad2a35dd02464c87a8645e23;
  assign mdsMatrix_54_6 = 253'h1bb04529d82ab5ee0345c9aa3132e3ffdc163696f871e9503f8a315052bef342;
  assign mdsMatrix_54_7 = 254'h344e8e15a9da104a0aeafbbf961dd2974015961b5c782d190d0b2918f2f4d6e7;
  assign mdsMatrix_54_8 = 252'h997ba24991e7b8b678b7ff0c755b98116856a56fa79deeaee122e076b536852;
  assign mdsMatrix_55_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_55_1 = 255'h514f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_55_2 = 255'h66d0f1e660ec4796f8b356e005810db9e6b5824adb6cc6dadb6db6dadb6db6dc;
  assign mdsMatrix_55_3 = 254'h2000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_55_4 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_55_5 = 251'h66269e6f2fa27dd10af9f8a1d64f50733cd4529556d65640000000eaaaaaa9c;
  assign mdsMatrix_55_6 = 254'h33321cd848c332c4bf155ed15280cc28ec9accfbb6a1c593b6db6d93b6db6dda;
  assign mdsMatrix_55_7 = 255'h40bb8a7ae0da4a8374247936b7210bdc6722d707495c966b4924926b49249227;
  assign mdsMatrix_55_8 = 255'h66369fb4d4c673ecf8389ab4f2f8bb12a0246b242c9cc9c9f3cf3ce665965973;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign tempAddrVec_5 = io_addr_regNext_5;
  assign tempAddrVec_6 = io_addr_regNext_6;
  assign tempAddrVec_7 = io_addr_regNext_7;
  assign tempAddrVec_8 = io_addr_regNext_8;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  assign io_data_5 = _zz_mdsMem_5_port0;
  assign io_data_6 = _zz_mdsMem_6_port0;
  assign io_data_7 = _zz_mdsMem_7_port0;
  assign io_data_8 = _zz_mdsMem_8_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
    io_addr_regNext_5 <= io_addr;
    io_addr_regNext_6 <= io_addr;
    io_addr_regNext_7 <= io_addr;
    io_addr_regNext_8 <= io_addr;
  end


endmodule

module MatrixConstantMem_8 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  input      [5:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire       [253:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [254:0]  mdsMatrix_0_2;
  wire       [254:0]  mdsMatrix_0_3;
  wire       [253:0]  mdsMatrix_0_4;
  wire       [253:0]  mdsMatrix_1_0;
  wire       [253:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [253:0]  mdsMatrix_1_3;
  wire       [254:0]  mdsMatrix_1_4;
  wire       [253:0]  mdsMatrix_2_0;
  wire       [253:0]  mdsMatrix_2_1;
  wire       [254:0]  mdsMatrix_2_2;
  wire       [253:0]  mdsMatrix_2_3;
  wire       [254:0]  mdsMatrix_2_4;
  wire       [253:0]  mdsMatrix_3_0;
  wire       [254:0]  mdsMatrix_3_1;
  wire       [253:0]  mdsMatrix_3_2;
  wire       [253:0]  mdsMatrix_3_3;
  wire       [254:0]  mdsMatrix_3_4;
  wire       [253:0]  mdsMatrix_4_0;
  wire       [252:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [254:0]  mdsMatrix_4_3;
  wire       [253:0]  mdsMatrix_4_4;
  wire       [253:0]  mdsMatrix_5_0;
  wire       [252:0]  mdsMatrix_5_1;
  wire       [251:0]  mdsMatrix_5_2;
  wire       [251:0]  mdsMatrix_5_3;
  wire       [252:0]  mdsMatrix_5_4;
  wire       [253:0]  mdsMatrix_6_0;
  wire       [254:0]  mdsMatrix_6_1;
  wire       [252:0]  mdsMatrix_6_2;
  wire       [254:0]  mdsMatrix_6_3;
  wire       [254:0]  mdsMatrix_6_4;
  wire       [253:0]  mdsMatrix_7_0;
  wire       [254:0]  mdsMatrix_7_1;
  wire       [254:0]  mdsMatrix_7_2;
  wire       [252:0]  mdsMatrix_7_3;
  wire       [254:0]  mdsMatrix_7_4;
  wire       [253:0]  mdsMatrix_8_0;
  wire       [253:0]  mdsMatrix_8_1;
  wire       [252:0]  mdsMatrix_8_2;
  wire       [253:0]  mdsMatrix_8_3;
  wire       [253:0]  mdsMatrix_8_4;
  wire       [253:0]  mdsMatrix_9_0;
  wire       [253:0]  mdsMatrix_9_1;
  wire       [254:0]  mdsMatrix_9_2;
  wire       [252:0]  mdsMatrix_9_3;
  wire       [253:0]  mdsMatrix_9_4;
  wire       [253:0]  mdsMatrix_10_0;
  wire       [253:0]  mdsMatrix_10_1;
  wire       [254:0]  mdsMatrix_10_2;
  wire       [252:0]  mdsMatrix_10_3;
  wire       [252:0]  mdsMatrix_10_4;
  wire       [253:0]  mdsMatrix_11_0;
  wire       [254:0]  mdsMatrix_11_1;
  wire       [247:0]  mdsMatrix_11_2;
  wire       [254:0]  mdsMatrix_11_3;
  wire       [254:0]  mdsMatrix_11_4;
  wire       [253:0]  mdsMatrix_12_0;
  wire       [254:0]  mdsMatrix_12_1;
  wire       [254:0]  mdsMatrix_12_2;
  wire       [251:0]  mdsMatrix_12_3;
  wire       [248:0]  mdsMatrix_12_4;
  wire       [253:0]  mdsMatrix_13_0;
  wire       [253:0]  mdsMatrix_13_1;
  wire       [253:0]  mdsMatrix_13_2;
  wire       [254:0]  mdsMatrix_13_3;
  wire       [252:0]  mdsMatrix_13_4;
  wire       [253:0]  mdsMatrix_14_0;
  wire       [253:0]  mdsMatrix_14_1;
  wire       [253:0]  mdsMatrix_14_2;
  wire       [253:0]  mdsMatrix_14_3;
  wire       [252:0]  mdsMatrix_14_4;
  wire       [253:0]  mdsMatrix_15_0;
  wire       [254:0]  mdsMatrix_15_1;
  wire       [251:0]  mdsMatrix_15_2;
  wire       [254:0]  mdsMatrix_15_3;
  wire       [251:0]  mdsMatrix_15_4;
  wire       [253:0]  mdsMatrix_16_0;
  wire       [253:0]  mdsMatrix_16_1;
  wire       [253:0]  mdsMatrix_16_2;
  wire       [254:0]  mdsMatrix_16_3;
  wire       [251:0]  mdsMatrix_16_4;
  wire       [253:0]  mdsMatrix_17_0;
  wire       [254:0]  mdsMatrix_17_1;
  wire       [250:0]  mdsMatrix_17_2;
  wire       [253:0]  mdsMatrix_17_3;
  wire       [252:0]  mdsMatrix_17_4;
  wire       [253:0]  mdsMatrix_18_0;
  wire       [253:0]  mdsMatrix_18_1;
  wire       [254:0]  mdsMatrix_18_2;
  wire       [253:0]  mdsMatrix_18_3;
  wire       [254:0]  mdsMatrix_18_4;
  wire       [253:0]  mdsMatrix_19_0;
  wire       [254:0]  mdsMatrix_19_1;
  wire       [252:0]  mdsMatrix_19_2;
  wire       [251:0]  mdsMatrix_19_3;
  wire       [254:0]  mdsMatrix_19_4;
  wire       [253:0]  mdsMatrix_20_0;
  wire       [254:0]  mdsMatrix_20_1;
  wire       [252:0]  mdsMatrix_20_2;
  wire       [252:0]  mdsMatrix_20_3;
  wire       [254:0]  mdsMatrix_20_4;
  wire       [253:0]  mdsMatrix_21_0;
  wire       [254:0]  mdsMatrix_21_1;
  wire       [252:0]  mdsMatrix_21_2;
  wire       [253:0]  mdsMatrix_21_3;
  wire       [253:0]  mdsMatrix_21_4;
  wire       [253:0]  mdsMatrix_22_0;
  wire       [253:0]  mdsMatrix_22_1;
  wire       [253:0]  mdsMatrix_22_2;
  wire       [252:0]  mdsMatrix_22_3;
  wire       [254:0]  mdsMatrix_22_4;
  wire       [253:0]  mdsMatrix_23_0;
  wire       [254:0]  mdsMatrix_23_1;
  wire       [252:0]  mdsMatrix_23_2;
  wire       [254:0]  mdsMatrix_23_3;
  wire       [254:0]  mdsMatrix_23_4;
  wire       [253:0]  mdsMatrix_24_0;
  wire       [254:0]  mdsMatrix_24_1;
  wire       [251:0]  mdsMatrix_24_2;
  wire       [252:0]  mdsMatrix_24_3;
  wire       [254:0]  mdsMatrix_24_4;
  wire       [253:0]  mdsMatrix_25_0;
  wire       [253:0]  mdsMatrix_25_1;
  wire       [252:0]  mdsMatrix_25_2;
  wire       [252:0]  mdsMatrix_25_3;
  wire       [254:0]  mdsMatrix_25_4;
  wire       [253:0]  mdsMatrix_26_0;
  wire       [254:0]  mdsMatrix_26_1;
  wire       [254:0]  mdsMatrix_26_2;
  wire       [248:0]  mdsMatrix_26_3;
  wire       [249:0]  mdsMatrix_26_4;
  wire       [253:0]  mdsMatrix_27_0;
  wire       [253:0]  mdsMatrix_27_1;
  wire       [254:0]  mdsMatrix_27_2;
  wire       [254:0]  mdsMatrix_27_3;
  wire       [252:0]  mdsMatrix_27_4;
  wire       [253:0]  mdsMatrix_28_0;
  wire       [254:0]  mdsMatrix_28_1;
  wire       [254:0]  mdsMatrix_28_2;
  wire       [250:0]  mdsMatrix_28_3;
  wire       [252:0]  mdsMatrix_28_4;
  wire       [253:0]  mdsMatrix_29_0;
  wire       [254:0]  mdsMatrix_29_1;
  wire       [253:0]  mdsMatrix_29_2;
  wire       [252:0]  mdsMatrix_29_3;
  wire       [253:0]  mdsMatrix_29_4;
  wire       [253:0]  mdsMatrix_30_0;
  wire       [252:0]  mdsMatrix_30_1;
  wire       [253:0]  mdsMatrix_30_2;
  wire       [254:0]  mdsMatrix_30_3;
  wire       [254:0]  mdsMatrix_30_4;
  wire       [253:0]  mdsMatrix_31_0;
  wire       [253:0]  mdsMatrix_31_1;
  wire       [254:0]  mdsMatrix_31_2;
  wire       [254:0]  mdsMatrix_31_3;
  wire       [253:0]  mdsMatrix_31_4;
  wire       [253:0]  mdsMatrix_32_0;
  wire       [254:0]  mdsMatrix_32_1;
  wire       [254:0]  mdsMatrix_32_2;
  wire       [254:0]  mdsMatrix_32_3;
  wire       [253:0]  mdsMatrix_32_4;
  wire       [253:0]  mdsMatrix_33_0;
  wire       [252:0]  mdsMatrix_33_1;
  wire       [253:0]  mdsMatrix_33_2;
  wire       [254:0]  mdsMatrix_33_3;
  wire       [253:0]  mdsMatrix_33_4;
  wire       [253:0]  mdsMatrix_34_0;
  wire       [254:0]  mdsMatrix_34_1;
  wire       [252:0]  mdsMatrix_34_2;
  wire       [254:0]  mdsMatrix_34_3;
  wire       [254:0]  mdsMatrix_34_4;
  wire       [253:0]  mdsMatrix_35_0;
  wire       [254:0]  mdsMatrix_35_1;
  wire       [253:0]  mdsMatrix_35_2;
  wire       [254:0]  mdsMatrix_35_3;
  wire       [252:0]  mdsMatrix_35_4;
  wire       [253:0]  mdsMatrix_36_0;
  wire       [252:0]  mdsMatrix_36_1;
  wire       [254:0]  mdsMatrix_36_2;
  wire       [254:0]  mdsMatrix_36_3;
  wire       [254:0]  mdsMatrix_36_4;
  wire       [253:0]  mdsMatrix_37_0;
  wire       [254:0]  mdsMatrix_37_1;
  wire       [250:0]  mdsMatrix_37_2;
  wire       [253:0]  mdsMatrix_37_3;
  wire       [252:0]  mdsMatrix_37_4;
  wire       [253:0]  mdsMatrix_38_0;
  wire       [253:0]  mdsMatrix_38_1;
  wire       [249:0]  mdsMatrix_38_2;
  wire       [254:0]  mdsMatrix_38_3;
  wire       [253:0]  mdsMatrix_38_4;
  wire       [253:0]  mdsMatrix_39_0;
  wire       [254:0]  mdsMatrix_39_1;
  wire       [252:0]  mdsMatrix_39_2;
  wire       [249:0]  mdsMatrix_39_3;
  wire       [253:0]  mdsMatrix_39_4;
  wire       [253:0]  mdsMatrix_40_0;
  wire       [250:0]  mdsMatrix_40_1;
  wire       [251:0]  mdsMatrix_40_2;
  wire       [254:0]  mdsMatrix_40_3;
  wire       [254:0]  mdsMatrix_40_4;
  wire       [253:0]  mdsMatrix_41_0;
  wire       [254:0]  mdsMatrix_41_1;
  wire       [253:0]  mdsMatrix_41_2;
  wire       [253:0]  mdsMatrix_41_3;
  wire       [252:0]  mdsMatrix_41_4;
  wire       [253:0]  mdsMatrix_42_0;
  wire       [254:0]  mdsMatrix_42_1;
  wire       [253:0]  mdsMatrix_42_2;
  wire       [253:0]  mdsMatrix_42_3;
  wire       [253:0]  mdsMatrix_42_4;
  wire       [253:0]  mdsMatrix_43_0;
  wire       [254:0]  mdsMatrix_43_1;
  wire       [254:0]  mdsMatrix_43_2;
  wire       [253:0]  mdsMatrix_43_3;
  wire       [254:0]  mdsMatrix_43_4;
  wire       [253:0]  mdsMatrix_44_0;
  wire       [253:0]  mdsMatrix_44_1;
  wire       [254:0]  mdsMatrix_44_2;
  wire       [253:0]  mdsMatrix_44_3;
  wire       [253:0]  mdsMatrix_44_4;
  wire       [253:0]  mdsMatrix_45_0;
  wire       [254:0]  mdsMatrix_45_1;
  wire       [248:0]  mdsMatrix_45_2;
  wire       [252:0]  mdsMatrix_45_3;
  wire       [254:0]  mdsMatrix_45_4;
  wire       [253:0]  mdsMatrix_46_0;
  wire       [254:0]  mdsMatrix_46_1;
  wire       [251:0]  mdsMatrix_46_2;
  wire       [253:0]  mdsMatrix_46_3;
  wire       [253:0]  mdsMatrix_46_4;
  wire       [253:0]  mdsMatrix_47_0;
  wire       [253:0]  mdsMatrix_47_1;
  wire       [253:0]  mdsMatrix_47_2;
  wire       [248:0]  mdsMatrix_47_3;
  wire       [254:0]  mdsMatrix_47_4;
  wire       [253:0]  mdsMatrix_48_0;
  wire       [248:0]  mdsMatrix_48_1;
  wire       [254:0]  mdsMatrix_48_2;
  wire       [251:0]  mdsMatrix_48_3;
  wire       [254:0]  mdsMatrix_48_4;
  wire       [253:0]  mdsMatrix_49_0;
  wire       [252:0]  mdsMatrix_49_1;
  wire       [253:0]  mdsMatrix_49_2;
  wire       [254:0]  mdsMatrix_49_3;
  wire       [252:0]  mdsMatrix_49_4;
  wire       [253:0]  mdsMatrix_50_0;
  wire       [253:0]  mdsMatrix_50_1;
  wire       [254:0]  mdsMatrix_50_2;
  wire       [253:0]  mdsMatrix_50_3;
  wire       [253:0]  mdsMatrix_50_4;
  wire       [253:0]  mdsMatrix_51_0;
  wire       [253:0]  mdsMatrix_51_1;
  wire       [254:0]  mdsMatrix_51_2;
  wire       [254:0]  mdsMatrix_51_3;
  wire       [252:0]  mdsMatrix_51_4;
  wire       [253:0]  mdsMatrix_52_0;
  wire       [252:0]  mdsMatrix_52_1;
  wire       [254:0]  mdsMatrix_52_2;
  wire       [250:0]  mdsMatrix_52_3;
  wire       [253:0]  mdsMatrix_52_4;
  wire       [253:0]  mdsMatrix_53_0;
  wire       [254:0]  mdsMatrix_53_1;
  wire       [246:0]  mdsMatrix_53_2;
  wire       [253:0]  mdsMatrix_53_3;
  wire       [254:0]  mdsMatrix_53_4;
  wire       [253:0]  mdsMatrix_54_0;
  wire       [254:0]  mdsMatrix_54_1;
  wire       [250:0]  mdsMatrix_54_2;
  wire       [254:0]  mdsMatrix_54_3;
  wire       [254:0]  mdsMatrix_54_4;
  wire       [5:0]    tempAddrVec_0;
  wire       [5:0]    tempAddrVec_1;
  wire       [5:0]    tempAddrVec_2;
  wire       [5:0]    tempAddrVec_3;
  wire       [5:0]    tempAddrVec_4;
  reg        [5:0]    io_addr_regNext;
  reg        [5:0]    io_addr_regNext_1;
  reg        [5:0]    io_addr_regNext_2;
  reg        [5:0]    io_addr_regNext_3;
  reg        [5:0]    io_addr_regNext_4;
  reg [254:0] mdsMem_0 [0:54];
  reg [254:0] mdsMem_1 [0:54];
  reg [254:0] mdsMem_2 [0:54];
  reg [254:0] mdsMem_3 [0:54];
  reg [254:0] mdsMem_4 [0:54];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_22_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_22_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_22_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_22_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_22_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  assign mdsMatrix_0_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_0_1 = 255'h653f541d0250843c3941db5d11e0dc68490f956aa21f233ecf63c74e844aa63d;
  assign mdsMatrix_0_2 = 255'h58d4574427df2005d4aba7f7f496a8c08bdabcd481f7fa79a8656ab26df5f222;
  assign mdsMatrix_0_3 = 255'h4f1a405f0b6791b3fc49ee7ca08ea2868510add04a5fd45d00228320ae8a1acd;
  assign mdsMatrix_0_4 = 254'h2a5e3dbd92b023b8c1ce42d02fb6daeccf3c6df3a88d490bcc321ecc11a9b553;
  assign mdsMatrix_1_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_1_1 = 254'h220e2bc9920aaab09a65d42a150beb75f47cb8b36072c059aef69cd2d0bc4304;
  assign mdsMatrix_1_2 = 255'h4fb8055ee30da4cc93eacd73c328b7cdcade8b9bf29e6a44a3fb8944b8ddfb65;
  assign mdsMatrix_1_3 = 254'h227985c374394938f17b36d606e4c9872bed2be3a26ed0e9ccb9ec2872a6d6c8;
  assign mdsMatrix_1_4 = 255'h583dc66284f5e1dd45c007374be177e61663e9bb1e60218a7eb7942819849847;
  assign mdsMatrix_2_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_2_1 = 254'h366a83c762e7da4da1c647842b246a09954a4946ca252264810fa97f1e46e652;
  assign mdsMatrix_2_2 = 255'h4579d0fea964e234bd8587f2ab211d81d587cd10b684ee6ee54e7b25c0147db5;
  assign mdsMatrix_2_3 = 254'h30a6da5372d92f633f57360b3af090d3b11f8933d036de7046991d41bd511123;
  assign mdsMatrix_2_4 = 255'h498e3f43f72255d7ac20d8a94d87380f44ae954831b1b4f121f011db3b5351ef;
  assign mdsMatrix_3_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_3_1 = 255'h49f4aaef6a1a7d2aaf5e352f88fdcb1b8bf2368e68cbaf88a4a2283fb90ad358;
  assign mdsMatrix_3_2 = 254'h3443a43b29202591730b46d31bda2edcb8386fc5d8b9ceebda682f163e02ceb4;
  assign mdsMatrix_3_3 = 254'h21951c4677852cd89d6980416678f7a4e1e99185a0dba0a4f1a4804b2fc03bc0;
  assign mdsMatrix_3_4 = 255'h682ec76748f8c5f6ed87108db463a11d346106c5ecd82d7d909d56a9898d393b;
  assign mdsMatrix_4_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_4_1 = 253'h11fa654f9df3670eee786b9eb8d37de4bd31db99e6ec7eae988daca33d4f0a24;
  assign mdsMatrix_4_2 = 255'h4a602ba9dbd595159790cf79d4dc3d1c696bba2e5faf3dfef189558a3fe21b15;
  assign mdsMatrix_4_3 = 255'h693ae8d0fcee12ba37ba806e972b27dcc5dd3bb547a423d7597f63d5429bd9c2;
  assign mdsMatrix_4_4 = 254'h3b1f83a3ef43909034dcbb2e0364884c184955fcb073b3bf618121c2e4c06778;
  assign mdsMatrix_5_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_5_1 = 253'h15805a671ec387f6c10ec5055eafadc08cf33b6cdfd8ab3620f536f3b418ea81;
  assign mdsMatrix_5_2 = 252'hc828efcdc38159fc39e17ad10c107a560957be3c354c03d9ef896af97bc56a3;
  assign mdsMatrix_5_3 = 252'hf7158dc2a3f7a118497b5adc82e795a4296a689b44565a8f77bcccb44838110;
  assign mdsMatrix_5_4 = 253'h1476d01de8d47f85884e25dbab81a83581fba6ce5c014c086c1564b33e10e3d6;
  assign mdsMatrix_6_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_6_1 = 255'h53ddbbd55b52f79f4670ab7e74db75849afdbf9928e3178cc47f075a2905d0f4;
  assign mdsMatrix_6_2 = 253'h1c5e70377e31a03c9837d055457d1f176082e508a79d1a35738d40e3a0f4eaae;
  assign mdsMatrix_6_3 = 255'h6af87023c24122c744082a23aad5d5ec630606fc447312de104f8689ed6161ec;
  assign mdsMatrix_6_4 = 255'h52c8653bd654fa155e01de602e00119a3d1d0273620aa85fbec8739026923c28;
  assign mdsMatrix_7_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_7_1 = 255'h6007092803a47e490dcfdc843a5b4e704b42ddad414d076f5f71f0f8cf2e6886;
  assign mdsMatrix_7_2 = 255'h568cdc2b19c623a84414310ff7abfe20a11b95f273c72ec98ed7d7c1ca519b7b;
  assign mdsMatrix_7_3 = 253'h13bbeedb5e9fca99411c5d7c7de1ffd957176beff35d46c5097594919c4dfb7a;
  assign mdsMatrix_7_4 = 255'h6af0a9153012462fd34cc300a97729fdef89abced0445e9fbc7308740e98ee40;
  assign mdsMatrix_8_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_8_1 = 254'h24d30f60b80b759777658e202a2b705b604ffd06f0b7b8efef0e71f1b5aff35a;
  assign mdsMatrix_8_2 = 253'h15e4110e1b7ea7c2e23396cf678dffb645eeca6066f8ed1a5100b6b734434f1a;
  assign mdsMatrix_8_3 = 254'h2cf4b1aef897d5cea96ad5dee203900a0e5b285b97a64163f6a227a7bb4b37df;
  assign mdsMatrix_8_4 = 254'h3ebab690698a00174ed67dbc7a0089077b4d877d895bbc5bd97344a25f2f08e7;
  assign mdsMatrix_9_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_9_1 = 254'h3c88b5e916b3bed6fe3edff2104fe45fcac40199c9176d2ea3923bbbe08037e3;
  assign mdsMatrix_9_2 = 255'h65ef3f0b5794773ab9febe6818ca6ce26042776fe632e101a2da63fc67ec3dd8;
  assign mdsMatrix_9_3 = 253'h1f09f4d47222fb924dbee66664a20d83ca7662412427d7cdde1a0ad61bb90420;
  assign mdsMatrix_9_4 = 254'h345628701ab9320b5bed04aa2de386d3a1bc95fd8e6b5aa9a9b19682146eaf28;
  assign mdsMatrix_10_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_10_1 = 254'h2758ab25e993e9a866cd0faa8ea70b8c5fb473678e26e5186babfab19a5c90c7;
  assign mdsMatrix_10_2 = 255'h6b5148e68b697f24511b0e6ad88d2df31d6a24b2a59409c921056cc7235f07fb;
  assign mdsMatrix_10_3 = 253'h16a8ba53c8b8e523f79e56dc0b59a79351908ceab008af56735e8a2f5e48846b;
  assign mdsMatrix_10_4 = 253'h1d36037010984f2a6a8cfcc90052a2167bab496c75cc997d741db5c869102bff;
  assign mdsMatrix_11_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_11_1 = 255'h50101f11a7e592689044447bb45b800eff12e3d61f0d35a89e7908ff8521408c;
  assign mdsMatrix_11_2 = 248'he37b374ada33eb17d0a22e0d870ecb7473ab0262db7c962e436ef8319d1734;
  assign mdsMatrix_11_3 = 255'h435d4ed58c8493436df63895cb6817793531e0d394b415505da064994f08aa5a;
  assign mdsMatrix_11_4 = 255'h57fec9efc6a769870c9f9d162d28f900f78eeea665052987424adba9edf603fa;
  assign mdsMatrix_12_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_12_1 = 255'h5179076cd15ea6437d4a295f206af51bea05c12abe05afd779c94c8ae884594e;
  assign mdsMatrix_12_2 = 255'h6861ecb95d0f7a41e9e8fc60c8ed06f87f09b263d64c5ef38b17da25a15be4e8;
  assign mdsMatrix_12_3 = 252'hcae818351438d4508bb99c2b77500536cfffa9afb60d4405981e365c8889a33;
  assign mdsMatrix_12_4 = 249'h1b771bc19961bf24d6bad9481f2477af19d2e6b398096702543e7014173d3d1;
  assign mdsMatrix_13_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_13_1 = 254'h304135ec1d9c7226d24239785798c917f1c2d8e4d0f2637a87f8de8e1fad04c7;
  assign mdsMatrix_13_2 = 254'h24c64c8a03fe4c3daba8d4c238a422123d4d884a1304d54a0459f36719e41215;
  assign mdsMatrix_13_3 = 255'h5bb368dfc57d231835ec58c5db5575dc75bca688801f018531b65c82bb8c7de1;
  assign mdsMatrix_13_4 = 253'h1b335bf96f73366229c73c251ad2b275f14b475a8d89c67c0e257190edd1fb02;
  assign mdsMatrix_14_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_14_1 = 254'h23c1e6343e79ce736c43210ad3bab1b51579940750841b780932d163089086aa;
  assign mdsMatrix_14_2 = 254'h3d2256c4f0e9531e19ad0ab8334b547aa4695d4f51df3a50be6508df8093e176;
  assign mdsMatrix_14_3 = 254'h2654a98c14f46d964bc71efba08e0dda0f31f6446469beb7b6f7834bc49cf636;
  assign mdsMatrix_14_4 = 253'h15edf1d71972352c288e5f942eb64aa98753485485006e096bd4812a7816efb2;
  assign mdsMatrix_15_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_15_1 = 255'h5a27495f68b2624243e7b244e6e0e7e28c896abb736999f248d9f2128c4fbcf4;
  assign mdsMatrix_15_2 = 252'hd9e20ead7ed2fc4dbe8104e400400c3fb9cdb488bce6f47dfc4f9098b037870;
  assign mdsMatrix_15_3 = 255'h589b4ad52cb5724d04dd9514a5c8d26d8d275dd97f94207afad4eb847f9aae87;
  assign mdsMatrix_15_4 = 252'hf0aa84c52408d8a6a322f640f9af2b09ff2969db6056abe64c183c368c81a84;
  assign mdsMatrix_16_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_16_1 = 254'h24266c14cb1c9fac578feca57f266021cbc27cf177a5a1d8a9a9eba99f380f3d;
  assign mdsMatrix_16_2 = 254'h21d3cc707395ff3794a6e4b6aa299bde3af22736f1b9697a831c91a7be018e9e;
  assign mdsMatrix_16_3 = 255'h520e8441933ec699c797cc21a05c928b85af0be0fc1da737cb7e095422737ca9;
  assign mdsMatrix_16_4 = 252'h8a2cf6b8a224f155b8f964804ca858ca24c6ec6c18d636cb832f0ef05c28e97;
  assign mdsMatrix_17_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_17_1 = 255'h62d83652f8c5d946d3a5d6b60aa4cb96e08d86c7d6536dd1be0a37a41623b94e;
  assign mdsMatrix_17_2 = 251'h58b5b09dd405514e66a43cce66bd2de42e6fbe9ccb230e5e2bc10026d8be376;
  assign mdsMatrix_17_3 = 254'h3c5b93f943baf3e774a0d559f133e0a43ae437604a256d58a543d4afc39563e6;
  assign mdsMatrix_17_4 = 253'h11ab86e56a37af61729ce74d095ae1686c698f9d64254abd60cd0b97c3846001;
  assign mdsMatrix_18_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_18_1 = 254'h31f50ccb2d5dff53301fad6d160480c93b19810bc967b774a0e9fdf0b45db37d;
  assign mdsMatrix_18_2 = 255'h73c6dc390861bbdad08661a4692a54849bbb0c2fade46b954cbe1d21ac65e6d4;
  assign mdsMatrix_18_3 = 254'h2a1105c95c28c093a55058f609616b4d17c95a58db408497757401cd47b3f0c8;
  assign mdsMatrix_18_4 = 255'h6ff3784e8d5eddda007b2e888107f8b4f35dc2b54b6baecd8ae58cb8366edb52;
  assign mdsMatrix_19_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_19_1 = 255'h61a44647a4bd8381651714023786737a5004f2bbf6b289033092a71a664ada81;
  assign mdsMatrix_19_2 = 253'h14460e2bdd0daebf92eafd4d6730b21d26effd60f6cd8dec8b325e52bf71fb85;
  assign mdsMatrix_19_3 = 252'hb9d5cc3e02da12fb3e9aff18d904cc6777c7a84eb9f11c9372c649d398bcc2d;
  assign mdsMatrix_19_4 = 255'h593fb4d01cdc0d79638f47c731e1aac21fb9cba453e25772fcc0515a6f27bb46;
  assign mdsMatrix_20_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_20_1 = 255'h6635475bf7e553adbfb4147c1a84e3b70829c94901a4f2a5f7cc1f20e1214f28;
  assign mdsMatrix_20_2 = 253'h16ac3a9d14d43af24f702a8d08b9d52131b482d193091bb62d47c5478acc599f;
  assign mdsMatrix_20_3 = 253'h18ed223e568da24d408635053ede53d0ef914de95f3ce510aca065f2b7a294d9;
  assign mdsMatrix_20_4 = 255'h53b0c9d77f358beeef457767f9c962b9e2ac5c47cba17d12e428f7d131d9ed8c;
  assign mdsMatrix_21_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_21_1 = 255'h48909ecd322c3966372bc3e516078d07b1a2420b8b41d5b616a60ee36fca233d;
  assign mdsMatrix_21_2 = 253'h10160d5d4275f05a276bd94bf3e5c35cb828ca0162c91aa74d34a8ebf3d54a3c;
  assign mdsMatrix_21_3 = 254'h22640b9956ba3ff4197aee826227e027585312b281c9021ff337f96ce03c4de5;
  assign mdsMatrix_21_4 = 254'h236e7b61b3b980df9d17a584e08776ef07074de269ea169db12cc6adca4c83e3;
  assign mdsMatrix_22_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_22_1 = 254'h3d8b71d044499381d88c722a4b5bdd9fae248e01e1da931d978fe6af9529e159;
  assign mdsMatrix_22_2 = 254'h3c1f49fd087dfb40f52e0fe3aa4d78fa4be7d1080155c8f06b9e115152242b67;
  assign mdsMatrix_22_3 = 253'h10a5cfa930afd11cc31e749f6c92e17426b1c0da9a8ae520a3819743c607bf29;
  assign mdsMatrix_22_4 = 255'h605c0f0f8ffd05badef96b0a12f912beec027b1bbd23416441d8de54e6d80772;
  assign mdsMatrix_23_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_23_1 = 255'h4b607b6b530075f5f0210d6bcfe4673ec1e958ebb539a3884983feb17fc6d824;
  assign mdsMatrix_23_2 = 253'h17c60d1040f80711e8d6f4d11be44100a7221a1d0b444a769b8dd0177f3fde4f;
  assign mdsMatrix_23_3 = 255'h5137c98c84baed98344e82c7fbe178c26ccd5f5c9c4b72526ff1434e5f258de0;
  assign mdsMatrix_23_4 = 255'h7125b032f6387fe1c06519cd5fe168761eb5eb2ae58888622ac0c528e0757c5b;
  assign mdsMatrix_24_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_24_1 = 255'h709b596a32f46aa53b6a01fa8c34ac125d05550d2ef9aad1167a61d0756b9c39;
  assign mdsMatrix_24_2 = 252'hfb82c92af10cadb3ab0b6121e1004ee421e383b6d65b29fd151e93171c18891;
  assign mdsMatrix_24_3 = 253'h178234f19d49b84de9abd5a749ed2506d6c57f32f8b71354260c1d4140f8f55e;
  assign mdsMatrix_24_4 = 255'h54e77827d33544c39e1eb11ded06a86493bb17f883fab9f6b73da761a9d3febf;
  assign mdsMatrix_25_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_25_1 = 254'h2a9ce0ea7c43212a6a96d4b86d97be6d68ce22cf4b0f1c7c18db7c953ee7d090;
  assign mdsMatrix_25_2 = 253'h15ada4802a9d66350d670fa4fa092702634e7fad2636cd239c3d4f01a83c48a4;
  assign mdsMatrix_25_3 = 253'h1e71fc25ad38700cbd24bbb850da52ac436ab65e9489f8dbfb7ba1bf5c7fca77;
  assign mdsMatrix_25_4 = 255'h57cffb79d22626dbb8ac73682e0caa0cb5e1cd64b6351fe169a94d8c049d1c87;
  assign mdsMatrix_26_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_26_1 = 255'h67ba354a3016c0f8bfa2cb86f8bff46db94915696dd668255008c9ae398b0e9e;
  assign mdsMatrix_26_2 = 255'h6c04b0e20df1932bf5ba10156521593eec23fcc30b59b522684d9315012e6b6f;
  assign mdsMatrix_26_3 = 249'h1672f634fccbb34bc11ea1b4970ab018cc6093ccd24b8d1bb5f9c353def7a0c;
  assign mdsMatrix_26_4 = 250'h3d15e99f8fc1b98eaaa28574fdc127339b9f15abefa355d5d94691589fafb27;
  assign mdsMatrix_27_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_27_1 = 254'h2c923f19105d15b62cbe727342bd304304cb228aeaf137dfb68b27227db2262d;
  assign mdsMatrix_27_2 = 255'h692a56b8ccd6103f7b380ee5c44886f96965c6f912b85771052757eff59fc37a;
  assign mdsMatrix_27_3 = 255'h59cb9986e1e54e5b62ee6c3c4e0ca039bb4f749d95a74130351241d1bcfbdbdf;
  assign mdsMatrix_27_4 = 253'h11572738860d65cd85238eb0a5370d3c25939cf90cb5d20b94376c17ff8ed09a;
  assign mdsMatrix_28_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_28_1 = 255'h515af7a94ee7a46ccb7d346480a82910d1b73ac9d59b661c1f9160eee4347e0a;
  assign mdsMatrix_28_2 = 255'h643e869950ed3e972cbdbb02f0443b7abba85980b4876a505494767dad211a9b;
  assign mdsMatrix_28_3 = 251'h5645bbb712c2988c5477f8ed487301d64d3797bd33ff91cc57349d8bf52b524;
  assign mdsMatrix_28_4 = 253'h1f3e7c40d6227fd9c1fcd885c43bb64fcd0825013f54218991d41a6950323029;
  assign mdsMatrix_29_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_29_1 = 255'h54a8537832b5ac47950cb00379ab564fd637cafe19d2b5a8d06ef4a86fc0cc1a;
  assign mdsMatrix_29_2 = 254'h3df1954b8e7479d31c3e0a4056f7cb8fcb8f084e7c45bc475ce320053986cc1a;
  assign mdsMatrix_29_3 = 253'h199b6d9c0586b27ee16436efeef329e0dde4dbeece6757cfb742f10988f6c5db;
  assign mdsMatrix_29_4 = 254'h20f6cef94174d57df374aaacd408a4bc3bf009ba19f7d06772b183e3b1706206;
  assign mdsMatrix_30_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_30_1 = 253'h1b8acd5cb580e6cbd4bc51117e30abc86cd2be0f3712743b5bb3c23862fc14e1;
  assign mdsMatrix_30_2 = 254'h225de8f2b850e57355f4bd1484629c73de1ad50a25ad25b1748ed2e5f4897c57;
  assign mdsMatrix_30_3 = 255'h675bad35f192cda3dc806ddbc13c14ea35182848a511fde4a6b381eb5290e294;
  assign mdsMatrix_30_4 = 255'h6410459755a2e1bb4c05accd16d3977b693ef6264494dc4f168c22a154bf475d;
  assign mdsMatrix_31_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_31_1 = 254'h3b206093ac93d859122ac618e1f9524adcfbb09bd0cffe16dd3b8eef0076aeea;
  assign mdsMatrix_31_2 = 255'h5e4d2914a520cb8f4d035f17e5f8d72583c26d39e975221583224833848d44fa;
  assign mdsMatrix_31_3 = 255'h670aa6a8784d7c24a29946ca276053933a8bdad2571b7a8fada1a84962e78603;
  assign mdsMatrix_31_4 = 254'h359a4cc6d4cdbbe86408da3d5c28979b340679e162429e5be20d5da5b23fa9dd;
  assign mdsMatrix_32_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_32_1 = 255'h71bc7ee2e44449a39b62ca673fc0e18776bdd4fd4fa5721dfbc14579979067c4;
  assign mdsMatrix_32_2 = 255'h6658d0ac36546fa37f5040115c1b6d7fb211800d854e42cc9ae3d30919b469c3;
  assign mdsMatrix_32_3 = 255'h4fc718c4bc7e90919cb9324735024bdbc1337e9dbb6538a31533a03264b061c8;
  assign mdsMatrix_32_4 = 254'h31ac4481291531ffeb397dd6d8d702a3a93ac6bdcd50caf418a90af2ecfeeb8e;
  assign mdsMatrix_33_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_33_1 = 253'h1708ec3065499a749eaa5aa39bcf58af5cc97b1fa612ad34f501bbfe7b8a33e3;
  assign mdsMatrix_33_2 = 254'h33f2de33a141a838a85787e3c4a9483ea5a71553e36c64dff3b8bf46f922fd1c;
  assign mdsMatrix_33_3 = 255'h5dca96e63cfb56d0f659dc6189dabbe406280340fae4fdf35daf0843086fe57c;
  assign mdsMatrix_33_4 = 254'h3583c9e97a514f391380bfb2f3b4f56831d35a42736b2e6e870e77b0e97ec43c;
  assign mdsMatrix_34_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_34_1 = 255'h4cd15bd787307b29464f0c0c7339e123a74fe02135d63d4b57ab467b7e78dadf;
  assign mdsMatrix_34_2 = 253'h16d7930f1b93251559607fc51aa97456b99981c8a3d5b349ee701362e7129713;
  assign mdsMatrix_34_3 = 255'h4a0c7a3a7e07593695cfa270480aa4e33c1937b2df0345ba293f04885bcda3f0;
  assign mdsMatrix_34_4 = 255'h4370a67fc9f798c063ee432ce20826f3dee702c63a4d3b9f96b79eaa28db9db6;
  assign mdsMatrix_35_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_35_1 = 255'h67e29d22eb037ecab605aea64002e4533432cbdc75d45aa10c7da8005fb9f6e9;
  assign mdsMatrix_35_2 = 254'h3a043f4ee071848a507bd6a31c39c7fee4418f511c0a8c9ecbd343b3b7292c20;
  assign mdsMatrix_35_3 = 255'h57e0d1b3bffebaeb16bce32ac1c03447ddd4f4244761fc25b26f7937192b98f1;
  assign mdsMatrix_35_4 = 253'h15f9caa21979edd55801987aa633b354e6cfdf0345e0e978df73f8f215232bc2;
  assign mdsMatrix_36_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_36_1 = 253'h17ddf3a806e30546c1c17955bf3b3a3f2473e5d1d9043f31950c970f0efb695c;
  assign mdsMatrix_36_2 = 255'h6bc5987764a24aa2847a2e29a555bbf77a8935bbf1c8b7f564e2d45ac5fae49d;
  assign mdsMatrix_36_3 = 255'h71fb1e5f5d00fe0c55cbc9014a27ffd3fc3a4823cd1e2b78c0655b54b3393f7c;
  assign mdsMatrix_36_4 = 255'h514533e8c085ed5ae95ddc9d0c8c3d33679cd938eb35a86c560ac3f45c8c4a69;
  assign mdsMatrix_37_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_37_1 = 255'h60932cdb234f4c4760bc9f1ed0d5eeb21fb8613d3f50aaf10ac8038120f68c85;
  assign mdsMatrix_37_2 = 251'h4205ea55d06ab113f67baa8b20f13d73d8100a0fd529ba20af51fbf98bc9c55;
  assign mdsMatrix_37_3 = 254'h207a1a3717b36742698bce4d5d66c73b51fd57d4d039b2c3d6f3eea8a233e5e6;
  assign mdsMatrix_37_4 = 253'h191622fc6c11e4c276574903fb6853c2cd3ba957191f0ebc07c949b112b5f6bc;
  assign mdsMatrix_38_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_38_1 = 254'h371b164d6eedcffd9772eed36e47bbb966a0e156b7dd7f1c978e6c2de2a28f3c;
  assign mdsMatrix_38_2 = 250'h33cdef197a30f3e46e34bfe364bcd36d2b5342d6c14a121f13860074f6a9f38;
  assign mdsMatrix_38_3 = 255'h6f25cf49f68d386c442970a82b54576cae60f7aa9cc27e78d6f477be5f4ad71b;
  assign mdsMatrix_38_4 = 254'h2a1e76206e844f96e7fd70a20b915282aa8767f9e956ba2f06762c351db4ee23;
  assign mdsMatrix_39_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_39_1 = 255'h50c62999c3da13f08781eba6074ffdbe78f406c99f52ce91afe54a9334d619f1;
  assign mdsMatrix_39_2 = 253'h1908f38263a4e682277a5fb87b917dd0a64b18aa9003c39820a9c931439b3c45;
  assign mdsMatrix_39_3 = 250'h2330d91dc2725fbd302e5d45dadfde601174fcb130b11cae7cd1f514b35a80b;
  assign mdsMatrix_39_4 = 254'h3c6c97f9f06d7880ff67aee054ff941424ad70fe049a03022ad81a457bbeb396;
  assign mdsMatrix_40_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_40_1 = 251'h7b9352af6d9c7cae2e3a8e4c451b31a76b748e9e3a60bf4e1f16567b132cc8a;
  assign mdsMatrix_40_2 = 252'hba9b61a620792c21cac8e4b19c3550e91e5a795113025e1dd0adf61352e0c96;
  assign mdsMatrix_40_3 = 255'h50114d3cfe233c2eeaf8d5439e25f7bd16713865d15f2a30e02ae881a3aa83cf;
  assign mdsMatrix_40_4 = 255'h590b5abe94890055ded5b5f9c0e20563bf3e14c83496b6b9d153583542c8c1db;
  assign mdsMatrix_41_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_41_1 = 255'h644a89d0c710fc3e02c8778f478898dd0fe43449f730ecdd8ad00f20f7f17e06;
  assign mdsMatrix_41_2 = 254'h29eb7427370a308be79f3debe74e8667a2911abf2d41877f3eaeb4abfda89a69;
  assign mdsMatrix_41_3 = 254'h2a7273922514078dd94191c90501b6fb3dcd8e13e5d6a78f0b7456cd5f105cce;
  assign mdsMatrix_41_4 = 253'h174e15da44ae13493995dcf7e67200584dd42d08ed74ab22b7130ec7e7ddab91;
  assign mdsMatrix_42_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_42_1 = 255'h5aecfbf6f9fbdf8e25799abf94af90c6f9e73641af2701b32efa6e67417df1c7;
  assign mdsMatrix_42_2 = 254'h341bc3e6ad146783eddeab8a6fc6b291c20cbc94c5c9c72ad54d6fe74dde9ecb;
  assign mdsMatrix_42_3 = 254'h3e9bf45493d4327b0f836c6611fb9bdcdfc0c8dc19cebb3b8fbc93d27dec7bf5;
  assign mdsMatrix_42_4 = 254'h2b86b3e7ae2aba18412ac4d3678e0d073fa16b7329c02a166b4cf8324f71a1e2;
  assign mdsMatrix_43_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_43_1 = 255'h5b26657c500fc2c0047345b31f5e7f617c0bfb9ae83349080e8fd50a2befbd38;
  assign mdsMatrix_43_2 = 255'h4134235dc375f5edd12fccc00472e5570764712d044b58f96ecb96c8edd3faca;
  assign mdsMatrix_43_3 = 254'h3a6b425bc8771fac301b181831aa9c8d067823f369fc06dc1d906910044ac4d7;
  assign mdsMatrix_43_4 = 255'h55a8691174f4ed92307b65a1b6001653af774f67aed54fc97c9e3c176362505c;
  assign mdsMatrix_44_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_44_1 = 254'h2fe05005372af070eda4a3b58aa706aca1fe55b8be6619245a201a6accad5195;
  assign mdsMatrix_44_2 = 255'h481b401ea1f4135b11eaa0d58cc184335ed26385bff24cd51e6bab5a1201a700;
  assign mdsMatrix_44_3 = 254'h296aceb16bcd1c8029992a074326a63bedf86606a144ac00abbfc9b1a27d34c3;
  assign mdsMatrix_44_4 = 254'h3455e45e6dc7b5be6580b8d4189c2b310b8166f51e72b6ebdfdf6f6d5e26b262;
  assign mdsMatrix_45_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_45_1 = 255'h5347ec0e340a13c5cd2c46422bbb586dc37826d96aa922836a4002fc24825efd;
  assign mdsMatrix_45_2 = 249'h1d5b922c9f98f44b016f5182f39977f8e9ccd4ac335da3e03a70153d3737780;
  assign mdsMatrix_45_3 = 253'h18bc0dc14cc3bd68d8629c03344eae503fa0b07fb66502c0fadca9d7d252b0d1;
  assign mdsMatrix_45_4 = 255'h5362639f9bf1cacf587f1be7577d1644ed6fd0939f39552d6745faaca26fbaa9;
  assign mdsMatrix_46_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_46_1 = 255'h723567d79678347acd0ddcc34e756bf09041d413dd8c5204b603030336f2c267;
  assign mdsMatrix_46_2 = 252'hed9af5906d3bfd0727eae2424f1a2951faf64f7a95358ab6fe2db1b32b7b709;
  assign mdsMatrix_46_3 = 254'h359f703813b1e4bc1eba428779cc9a949a3877441ce188366584988be7454b02;
  assign mdsMatrix_46_4 = 254'h235b1a204e94453b20dcfef2291b7b181c0138127e4983943277eac8a7f92bf2;
  assign mdsMatrix_47_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_47_1 = 254'h31bb21d3d08a250c3defcaf73783f3b25f4a310ce14107443206628907fc8a74;
  assign mdsMatrix_47_2 = 254'h2deecea2bc7e68cf83df00dc972c2b19194a898befd0e435d4d73573d9b4b50d;
  assign mdsMatrix_47_3 = 249'h128fbf471e30672a6ed09ed0cdc303aa0e124ee2be43e81942e815fb0a6520f;
  assign mdsMatrix_47_4 = 255'h60cb3eb713da2e123a98b16fad3e335cf7fec1cd16d995e09208c10eb259cfbc;
  assign mdsMatrix_48_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_48_1 = 249'h1403362fb2102129307110f40570ef437778055a8540fc493f36f4b0754d4ec;
  assign mdsMatrix_48_2 = 255'h5836c684049360b133c7c210ee8bec32c8d865144a5773157a9bc9aac0b8a59b;
  assign mdsMatrix_48_3 = 252'h8a2c2c1530b892638cd889f5a897b4588313ee2aeb86c25cf934b1e2ffd085e;
  assign mdsMatrix_48_4 = 255'h6ea0c47c01a3ad02a436aa75047167f6eba4e778416e6c7dfccc0c9136eb9912;
  assign mdsMatrix_49_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_49_1 = 253'h10e28ea08183764284ce21cb80521557ed8e8b6f5e5b75fb735ed211102ddd68;
  assign mdsMatrix_49_2 = 254'h38ccba5cc6b9fce48b228c38edd5c1b961fa237e1a566ea053a93946b22c5a3f;
  assign mdsMatrix_49_3 = 255'h70e867288781fa5b71d7f5a0342756cc635f2dd4d882c6a44b1d5561b4e267fd;
  assign mdsMatrix_49_4 = 253'h1c48ba2daa6b59fb569119077842b7f883629698c4f1673cc6b5b2e2d2e435bd;
  assign mdsMatrix_50_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_50_1 = 254'h25d6bcc3903c6202a6feb6ce060c115ad91341c3bce9e0fb7ddab7b437dda5bf;
  assign mdsMatrix_50_2 = 255'h664651c66ca4e8759c20ac3764eb8e717b259db286a50de9b6cc0ff41e093658;
  assign mdsMatrix_50_3 = 254'h3e12f6eceea7ef2fb490761b29e5ac8fa0c2c267106407bbc135376c3ecac86c;
  assign mdsMatrix_50_4 = 254'h2fb3498cd03a8e6118082a0b34513ea83b5ef727a7d66823d9ab094ef321c3ad;
  assign mdsMatrix_51_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_51_1 = 254'h3833a6fdf04f6034c1fd6f683e8b856e27c33eab603c6a9d8a6413f7a449f69b;
  assign mdsMatrix_51_2 = 255'h5a08a632c1ac8d7215a574b8a03fe0001ae44360939a285bb3750310bd3f8759;
  assign mdsMatrix_51_3 = 255'h560ebe981d37ca4b2b8bd4c7968ea75dea912d0352728b4d17b8374ce847c8b3;
  assign mdsMatrix_51_4 = 253'h16ae2f7053b1f2ee97c6aa12b37ca3ceb374026020cdb305e3de416c828824fa;
  assign mdsMatrix_52_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_52_1 = 253'h13c6c19a7304cef1d9a4b83b61c032f2c2557c2a95892b401861861845e45e46;
  assign mdsMatrix_52_2 = 255'h68ced4716687cdcb90f6074ef0a191ce6ea455655ac8d9662116a3b285dcf019;
  assign mdsMatrix_52_3 = 251'h588d372db0b48c6c5d77f6e3abddbb485ec6aff38174708000e2707fff1d8f8;
  assign mdsMatrix_52_4 = 254'h2a6cbe351fd6c0ca4664a70116525b7d8fa0a4e443301feeffef37223343fc11;
  assign mdsMatrix_53_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_53_1 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_53_2 = 247'h50d08f5d9edbd7bdae0af775ffb812b1693296b46b86b49249249270270270;
  assign mdsMatrix_53_3 = 254'h233a465de57dff1e94962bfe80a642ed79764e9e0de1a07600000875fffff78a;
  assign mdsMatrix_53_4 = 255'h43b51c27d123d0e9f0877396bcb0f21456b3f93455fdb465fffff5ff9999a39a;
  assign mdsMatrix_54_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_54_1 = 255'h4000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_54_2 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_54_3 = 255'h486e140d064f104ecca4efcfc634efe0098e27ee0009d80600000005fffffffa;
  assign mdsMatrix_54_4 = 255'h413a32e3a532f1ddd72cc9c36549968219da21a9332aab2dfffffffaccccccd2;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
  end


endmodule

module MatrixConstantMem_7 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  output     [254:0]  io_data_9,
  output     [254:0]  io_data_10,
  output     [254:0]  io_data_11,
  input      [3:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  reg        [254:0]  _zz_mdsMem_5_port0;
  reg        [254:0]  _zz_mdsMem_6_port0;
  reg        [254:0]  _zz_mdsMem_7_port0;
  reg        [254:0]  _zz_mdsMem_8_port0;
  reg        [254:0]  _zz_mdsMem_9_port0;
  reg        [254:0]  _zz_mdsMem_10_port0;
  reg        [254:0]  _zz_mdsMem_11_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire                _zz_mdsMem_5_port;
  wire                _zz_io_data_5;
  wire                _zz_mdsMem_6_port;
  wire                _zz_io_data_6;
  wire                _zz_mdsMem_7_port;
  wire                _zz_io_data_7;
  wire                _zz_mdsMem_8_port;
  wire                _zz_io_data_8;
  wire                _zz_mdsMem_9_port;
  wire                _zz_io_data_9;
  wire                _zz_mdsMem_10_port;
  wire                _zz_io_data_10;
  wire                _zz_mdsMem_11_port;
  wire                _zz_io_data_11;
  wire       [254:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [252:0]  mdsMatrix_0_2;
  wire       [250:0]  mdsMatrix_0_3;
  wire       [253:0]  mdsMatrix_0_4;
  wire       [254:0]  mdsMatrix_0_5;
  wire       [250:0]  mdsMatrix_0_6;
  wire       [254:0]  mdsMatrix_0_7;
  wire       [254:0]  mdsMatrix_0_8;
  wire       [254:0]  mdsMatrix_0_9;
  wire       [254:0]  mdsMatrix_0_10;
  wire       [254:0]  mdsMatrix_0_11;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [252:0]  mdsMatrix_1_1;
  wire       [253:0]  mdsMatrix_1_2;
  wire       [253:0]  mdsMatrix_1_3;
  wire       [253:0]  mdsMatrix_1_4;
  wire       [253:0]  mdsMatrix_1_5;
  wire       [252:0]  mdsMatrix_1_6;
  wire       [254:0]  mdsMatrix_1_7;
  wire       [254:0]  mdsMatrix_1_8;
  wire       [253:0]  mdsMatrix_1_9;
  wire       [252:0]  mdsMatrix_1_10;
  wire       [254:0]  mdsMatrix_1_11;
  wire       [253:0]  mdsMatrix_2_0;
  wire       [253:0]  mdsMatrix_2_1;
  wire       [252:0]  mdsMatrix_2_2;
  wire       [253:0]  mdsMatrix_2_3;
  wire       [254:0]  mdsMatrix_2_4;
  wire       [254:0]  mdsMatrix_2_5;
  wire       [253:0]  mdsMatrix_2_6;
  wire       [254:0]  mdsMatrix_2_7;
  wire       [253:0]  mdsMatrix_2_8;
  wire       [253:0]  mdsMatrix_2_9;
  wire       [254:0]  mdsMatrix_2_10;
  wire       [253:0]  mdsMatrix_2_11;
  wire       [254:0]  mdsMatrix_3_0;
  wire       [253:0]  mdsMatrix_3_1;
  wire       [253:0]  mdsMatrix_3_2;
  wire       [253:0]  mdsMatrix_3_3;
  wire       [252:0]  mdsMatrix_3_4;
  wire       [253:0]  mdsMatrix_3_5;
  wire       [253:0]  mdsMatrix_3_6;
  wire       [254:0]  mdsMatrix_3_7;
  wire       [254:0]  mdsMatrix_3_8;
  wire       [254:0]  mdsMatrix_3_9;
  wire       [252:0]  mdsMatrix_3_10;
  wire       [254:0]  mdsMatrix_3_11;
  wire       [252:0]  mdsMatrix_4_0;
  wire       [253:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [252:0]  mdsMatrix_4_3;
  wire       [253:0]  mdsMatrix_4_4;
  wire       [254:0]  mdsMatrix_4_5;
  wire       [252:0]  mdsMatrix_4_6;
  wire       [253:0]  mdsMatrix_4_7;
  wire       [254:0]  mdsMatrix_4_8;
  wire       [253:0]  mdsMatrix_4_9;
  wire       [252:0]  mdsMatrix_4_10;
  wire       [254:0]  mdsMatrix_4_11;
  wire       [253:0]  mdsMatrix_5_0;
  wire       [253:0]  mdsMatrix_5_1;
  wire       [254:0]  mdsMatrix_5_2;
  wire       [253:0]  mdsMatrix_5_3;
  wire       [254:0]  mdsMatrix_5_4;
  wire       [252:0]  mdsMatrix_5_5;
  wire       [253:0]  mdsMatrix_5_6;
  wire       [252:0]  mdsMatrix_5_7;
  wire       [252:0]  mdsMatrix_5_8;
  wire       [254:0]  mdsMatrix_5_9;
  wire       [253:0]  mdsMatrix_5_10;
  wire       [253:0]  mdsMatrix_5_11;
  wire       [254:0]  mdsMatrix_6_0;
  wire       [252:0]  mdsMatrix_6_1;
  wire       [253:0]  mdsMatrix_6_2;
  wire       [253:0]  mdsMatrix_6_3;
  wire       [252:0]  mdsMatrix_6_4;
  wire       [253:0]  mdsMatrix_6_5;
  wire       [252:0]  mdsMatrix_6_6;
  wire       [253:0]  mdsMatrix_6_7;
  wire       [253:0]  mdsMatrix_6_8;
  wire       [253:0]  mdsMatrix_6_9;
  wire       [254:0]  mdsMatrix_6_10;
  wire       [254:0]  mdsMatrix_6_11;
  wire       [252:0]  mdsMatrix_7_0;
  wire       [254:0]  mdsMatrix_7_1;
  wire       [254:0]  mdsMatrix_7_2;
  wire       [254:0]  mdsMatrix_7_3;
  wire       [253:0]  mdsMatrix_7_4;
  wire       [252:0]  mdsMatrix_7_5;
  wire       [253:0]  mdsMatrix_7_6;
  wire       [253:0]  mdsMatrix_7_7;
  wire       [252:0]  mdsMatrix_7_8;
  wire       [254:0]  mdsMatrix_7_9;
  wire       [254:0]  mdsMatrix_7_10;
  wire       [254:0]  mdsMatrix_7_11;
  wire       [253:0]  mdsMatrix_8_0;
  wire       [254:0]  mdsMatrix_8_1;
  wire       [253:0]  mdsMatrix_8_2;
  wire       [254:0]  mdsMatrix_8_3;
  wire       [254:0]  mdsMatrix_8_4;
  wire       [252:0]  mdsMatrix_8_5;
  wire       [253:0]  mdsMatrix_8_6;
  wire       [252:0]  mdsMatrix_8_7;
  wire       [254:0]  mdsMatrix_8_8;
  wire       [254:0]  mdsMatrix_8_9;
  wire       [254:0]  mdsMatrix_8_10;
  wire       [253:0]  mdsMatrix_8_11;
  wire       [254:0]  mdsMatrix_9_0;
  wire       [253:0]  mdsMatrix_9_1;
  wire       [253:0]  mdsMatrix_9_2;
  wire       [254:0]  mdsMatrix_9_3;
  wire       [253:0]  mdsMatrix_9_4;
  wire       [254:0]  mdsMatrix_9_5;
  wire       [253:0]  mdsMatrix_9_6;
  wire       [254:0]  mdsMatrix_9_7;
  wire       [254:0]  mdsMatrix_9_8;
  wire       [254:0]  mdsMatrix_9_9;
  wire       [252:0]  mdsMatrix_9_10;
  wire       [253:0]  mdsMatrix_9_11;
  wire       [252:0]  mdsMatrix_10_0;
  wire       [252:0]  mdsMatrix_10_1;
  wire       [254:0]  mdsMatrix_10_2;
  wire       [252:0]  mdsMatrix_10_3;
  wire       [252:0]  mdsMatrix_10_4;
  wire       [253:0]  mdsMatrix_10_5;
  wire       [254:0]  mdsMatrix_10_6;
  wire       [254:0]  mdsMatrix_10_7;
  wire       [254:0]  mdsMatrix_10_8;
  wire       [252:0]  mdsMatrix_10_9;
  wire       [254:0]  mdsMatrix_10_10;
  wire       [254:0]  mdsMatrix_10_11;
  wire       [250:0]  mdsMatrix_11_0;
  wire       [254:0]  mdsMatrix_11_1;
  wire       [253:0]  mdsMatrix_11_2;
  wire       [254:0]  mdsMatrix_11_3;
  wire       [254:0]  mdsMatrix_11_4;
  wire       [253:0]  mdsMatrix_11_5;
  wire       [254:0]  mdsMatrix_11_6;
  wire       [254:0]  mdsMatrix_11_7;
  wire       [253:0]  mdsMatrix_11_8;
  wire       [253:0]  mdsMatrix_11_9;
  wire       [254:0]  mdsMatrix_11_10;
  wire       [254:0]  mdsMatrix_11_11;
  wire       [3:0]    tempAddrVec_0;
  wire       [3:0]    tempAddrVec_1;
  wire       [3:0]    tempAddrVec_2;
  wire       [3:0]    tempAddrVec_3;
  wire       [3:0]    tempAddrVec_4;
  wire       [3:0]    tempAddrVec_5;
  wire       [3:0]    tempAddrVec_6;
  wire       [3:0]    tempAddrVec_7;
  wire       [3:0]    tempAddrVec_8;
  wire       [3:0]    tempAddrVec_9;
  wire       [3:0]    tempAddrVec_10;
  wire       [3:0]    tempAddrVec_11;
  reg        [3:0]    io_addr_regNext;
  reg        [3:0]    io_addr_regNext_1;
  reg        [3:0]    io_addr_regNext_2;
  reg        [3:0]    io_addr_regNext_3;
  reg        [3:0]    io_addr_regNext_4;
  reg        [3:0]    io_addr_regNext_5;
  reg        [3:0]    io_addr_regNext_6;
  reg        [3:0]    io_addr_regNext_7;
  reg        [3:0]    io_addr_regNext_8;
  reg        [3:0]    io_addr_regNext_9;
  reg        [3:0]    io_addr_regNext_10;
  reg        [3:0]    io_addr_regNext_11;
  reg [254:0] mdsMem_0 [0:11];
  reg [254:0] mdsMem_1 [0:11];
  reg [254:0] mdsMem_2 [0:11];
  reg [254:0] mdsMem_3 [0:11];
  reg [254:0] mdsMem_4 [0:11];
  reg [254:0] mdsMem_5 [0:11];
  reg [254:0] mdsMem_6 [0:11];
  reg [254:0] mdsMem_7 [0:11];
  reg [254:0] mdsMem_8 [0:11];
  reg [254:0] mdsMem_9 [0:11];
  reg [254:0] mdsMem_10 [0:11];
  reg [254:0] mdsMem_11 [0:11];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  assign _zz_io_data_5 = 1'b1;
  assign _zz_io_data_6 = 1'b1;
  assign _zz_io_data_7 = 1'b1;
  assign _zz_io_data_8 = 1'b1;
  assign _zz_io_data_9 = 1'b1;
  assign _zz_io_data_10 = 1'b1;
  assign _zz_io_data_11 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_5.bin",mdsMem_5);
  end
  always @(posedge clk) begin
    if(_zz_io_data_5) begin
      _zz_mdsMem_5_port0 <= mdsMem_5[tempAddrVec_5];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_6.bin",mdsMem_6);
  end
  always @(posedge clk) begin
    if(_zz_io_data_6) begin
      _zz_mdsMem_6_port0 <= mdsMem_6[tempAddrVec_6];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_7.bin",mdsMem_7);
  end
  always @(posedge clk) begin
    if(_zz_io_data_7) begin
      _zz_mdsMem_7_port0 <= mdsMem_7[tempAddrVec_7];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_8.bin",mdsMem_8);
  end
  always @(posedge clk) begin
    if(_zz_io_data_8) begin
      _zz_mdsMem_8_port0 <= mdsMem_8[tempAddrVec_8];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_9.bin",mdsMem_9);
  end
  always @(posedge clk) begin
    if(_zz_io_data_9) begin
      _zz_mdsMem_9_port0 <= mdsMem_9[tempAddrVec_9];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_10.bin",mdsMem_10);
  end
  always @(posedge clk) begin
    if(_zz_io_data_10) begin
      _zz_mdsMem_10_port0 <= mdsMem_10[tempAddrVec_10];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_21_mdsMem_11.bin",mdsMem_11);
  end
  always @(posedge clk) begin
    if(_zz_io_data_11) begin
      _zz_mdsMem_11_port0 <= mdsMem_11[tempAddrVec_11];
    end
  end

  assign mdsMatrix_0_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_0_1 = 255'h47c5564e1a68586b0a8728b66a7179dab86caac297ff58013b3d2a20f1c99be7;
  assign mdsMatrix_0_2 = 253'h163b11236936498bb83f8693199c1b42bdc4c2a16ad0cf319328fb56f5fff37c;
  assign mdsMatrix_0_3 = 251'h67e187f6bab44d5464d50f593bb130b15080a0c3f862a16cfe8be4c1c09eb2f;
  assign mdsMatrix_0_4 = 254'h3bc66b1bb15314767aba0afe5e2a415458351e9ecbb7703b3799e2a277874120;
  assign mdsMatrix_0_5 = 255'h616800830f8f6c24350a0742a1cde0ac8f1ceadea689604a2944831325861aaa;
  assign mdsMatrix_0_6 = 251'h45eb10a19acbd075876279c36e6655e3cdf5f55a719c84b04265e0646fc0353;
  assign mdsMatrix_0_7 = 255'h4192893c761c0a4bd6d8e66cb23779bafc4e7b9b320cbe6a079da190acdc8167;
  assign mdsMatrix_0_8 = 255'h673373d1c03971e7e5aefee9e711cbae205847c251d669f4845a659feb773e40;
  assign mdsMatrix_0_9 = 255'h6d4072b155434516531282095c6f4947204b5601e1b43a623e5b6f07e2cdc6bc;
  assign mdsMatrix_0_10 = 255'h5ca95e2061b8f68927f732b4966ca50cf88ea7ccf27298ec3c43fac1ec031c0b;
  assign mdsMatrix_0_11 = 255'h6689c92e2cb339add91b4cabe6e59144daf07e94e173351fbff5ed22317d0efb;
  assign mdsMatrix_1_0 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_1_1 = 253'h15c7927460f1e76ade9fac71e5ce4acdc964f5ffadd55b14f465d9696dc20d1b;
  assign mdsMatrix_1_2 = 254'h2d99595949d2bb6dec34d0ae1be5305aecbea2ac862370cafcb805f20f6329ca;
  assign mdsMatrix_1_3 = 254'h34829997b5e1d50eef6933882583126ac9fec1f5734c5bd50fe3fbf12a8b9c8f;
  assign mdsMatrix_1_4 = 254'h314863966fb120a682b548e166e07a305b0dd5ab573bdaecc5a5cde6107c23e9;
  assign mdsMatrix_1_5 = 254'h3f6474544054fdd06fc462d66a0ba8fd31aafcc5fc7baa4abb9db3519aff0eb8;
  assign mdsMatrix_1_6 = 253'h158b2694a1ea2cd8a80374af820c8dbc9711bc56537ee77c8012960c9d2842bb;
  assign mdsMatrix_1_7 = 255'h5926065232ef9bedc453194039fc15e36da21887af005004ee3fd2cc28aef675;
  assign mdsMatrix_1_8 = 255'h72a1062b57f4fa2e5771859d22f5fcd86130db83e0d506225b103cc5d3074aa7;
  assign mdsMatrix_1_9 = 254'h31d6995c6cfbe12818215b4349112482433988d1570f2c621c9e671a7684a3ef;
  assign mdsMatrix_1_10 = 253'h14ff39ce71663ed6904498dc2b0cd2ffdd9f3da50d3b747d587adbd1ff4e192d;
  assign mdsMatrix_1_11 = 255'h6a758500fad34882feffcb009873e6077e78d4300020f33ef22f40faba7981f7;
  assign mdsMatrix_2_0 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_2_1 = 254'h2d99595949d2bb6dec34d0ae1be5305aecbea2ac862370cafcb805f20f6329ca;
  assign mdsMatrix_2_2 = 253'h10b3b3bfab132caad43f673a621a415b26bcd16e5815d48dfb6d736099db78cb;
  assign mdsMatrix_2_3 = 254'h2ef0f7816ba3fac16753784ff247aa251fa6cab899dba1fd792d5cf8821c8854;
  assign mdsMatrix_2_4 = 255'h654416d02749658d519a50a707c0fc5b2de6fcb167b3b45726c48c22eae61fdd;
  assign mdsMatrix_2_5 = 255'h660387e933bce0aa3c0a7ed289144f5f6409672e58703eb83e4676c83710b1bd;
  assign mdsMatrix_2_6 = 254'h30094b90300c289449619e9be98b827b619d4d7e8ddc460362949e9daeca7116;
  assign mdsMatrix_2_7 = 255'h41ee23f17d0025d61cd2578b9b47d8e2034c1999863c94b2b086e23a0c695685;
  assign mdsMatrix_2_8 = 254'h3cc52207bbd8577c030f4eb9521656c95a079c6c229005a7d5641c2e65c04144;
  assign mdsMatrix_2_9 = 254'h29ff2b59e1bc0353ecaf1d87cc085f91c8ed9b6212448aa1b5ceec55c996d003;
  assign mdsMatrix_2_10 = 255'h5270a6310562c5907877e43b1bfa6e064ffdc02a8ec763fcf472d48e39acbd42;
  assign mdsMatrix_2_11 = 254'h349cdd4bc00a305e5677872bbed238d65beae70b5f35522b3642560b63a5d7f0;
  assign mdsMatrix_3_0 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_3_1 = 254'h34829997b5e1d50eef6933882583126ac9fec1f5734c5bd50fe3fbf12a8b9c8f;
  assign mdsMatrix_3_2 = 254'h2ef0f7816ba3fac16753784ff247aa251fa6cab899dba1fd792d5cf8821c8854;
  assign mdsMatrix_3_3 = 254'h21f3df4240ce99eb77f4a8b1c5d1be9ae815e4507f73d63851eb8f798362e97e;
  assign mdsMatrix_3_4 = 253'h17bfd17b0aad4c6c59d072382da3b36d6adf091531e6b10cd8159289c0f23c34;
  assign mdsMatrix_3_5 = 254'h25c7568d870c388fa5fd85d9a44bf5935f49f677f2da648e10f82bf27ee4b644;
  assign mdsMatrix_3_6 = 254'h2ad34bcfe341c5685c018acf0b5a7c11d9649534ca1e6c65c7432b4b0e646874;
  assign mdsMatrix_3_7 = 255'h69d9f9f632557ac2c4ce207d2a80dc053bd63a7d505b1a8f93281484f38af5ba;
  assign mdsMatrix_3_8 = 255'h4177ffe5b5c4a55c525b37d5ec1f55eda6fade24205b20ba52cba1d4eb3d52b9;
  assign mdsMatrix_3_9 = 255'h67e14645d098f70fa8c0e28a73bd0f75eceb766df2373013b1781684b482c9fb;
  assign mdsMatrix_3_10 = 253'h197ba23e784e407b5d5513b59adbb98fa16dcb92bb6943197d3760b49b1dd1d1;
  assign mdsMatrix_3_11 = 255'h5753b589f9a06db49d750abe1351345af62a29ee5b6714168fc9785e6be004d3;
  assign mdsMatrix_4_0 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_4_1 = 254'h314863966fb120a682b548e166e07a305b0dd5ab573bdaecc5a5cde6107c23e9;
  assign mdsMatrix_4_2 = 255'h654416d02749658d519a50a707c0fc5b2de6fcb167b3b45726c48c22eae61fdd;
  assign mdsMatrix_4_3 = 253'h17bfd17b0aad4c6c59d072382da3b36d6adf091531e6b10cd8159289c0f23c34;
  assign mdsMatrix_4_4 = 254'h2eb096014ec9c7774548a5f6e1326cce03ca54b5fbea384d6546534ab395e095;
  assign mdsMatrix_4_5 = 255'h59a0690d52f046fa0382894b468794aa857a9ce17d25589e1cc541a7813d0e2e;
  assign mdsMatrix_4_6 = 253'h173346c563ec6dbe554f8b0221dbfc5da410af5cce0f15e4949f788f1c24cfde;
  assign mdsMatrix_4_7 = 254'h251e29d5bcec361c6a65da991cfb90f96f9f7c650bd94876f09fe8c9ab2c354c;
  assign mdsMatrix_4_8 = 255'h4ebf8c6b40211b8a277d5a9d9d1014c18582596cf8ac3812e752af8428ba98e0;
  assign mdsMatrix_4_9 = 254'h3ccfb0b82d30e2a96b4c21ed0cffffc34673eda2395e1b8db9cde8ab0e59d519;
  assign mdsMatrix_4_10 = 253'h1ee8136953d9562ca3d0eb11698492c3c038b41c27d30886b5f4111f8a4e6c68;
  assign mdsMatrix_4_11 = 255'h73a64e645c8c1cd18133f48ab3afdb4d1fae4241e83c6a4d429aa513f9a3414b;
  assign mdsMatrix_5_0 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_5_1 = 254'h3f6474544054fdd06fc462d66a0ba8fd31aafcc5fc7baa4abb9db3519aff0eb8;
  assign mdsMatrix_5_2 = 255'h660387e933bce0aa3c0a7ed289144f5f6409672e58703eb83e4676c83710b1bd;
  assign mdsMatrix_5_3 = 254'h25c7568d870c388fa5fd85d9a44bf5935f49f677f2da648e10f82bf27ee4b644;
  assign mdsMatrix_5_4 = 255'h59a0690d52f046fa0382894b468794aa857a9ce17d25589e1cc541a7813d0e2e;
  assign mdsMatrix_5_5 = 253'h119047bef9dded3e553eb68845d89e887afba808ab64fb0213288e785c4c67d0;
  assign mdsMatrix_5_6 = 254'h284b46d9e6433e109fa41b53ef70ce50a47c184a41bda636d92727ec0fa535f8;
  assign mdsMatrix_5_7 = 253'h15064f004897e03209e30a2f225c50005d634ee8086ab971be720ed7339b8180;
  assign mdsMatrix_5_8 = 253'h1ae7d0b1501894960d8ef684c43bb9392c60c9f7c465d26081631de66ab866ef;
  assign mdsMatrix_5_9 = 255'h4f6b915cd211c03922929e2bcda92d5d62c827224dbb0ec3ca13da4488dad173;
  assign mdsMatrix_5_10 = 254'h2f9e31da3bca17f740ab3b2e13254875e6337da40fd7e6b76bfc9d776809c972;
  assign mdsMatrix_5_11 = 254'h39480b0425cd85cec7d8f43d000238cc3ca6805ba6fe7d8248330dc9bcdd1f18;
  assign mdsMatrix_6_0 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_6_1 = 253'h158b2694a1ea2cd8a80374af820c8dbc9711bc56537ee77c8012960c9d2842bb;
  assign mdsMatrix_6_2 = 254'h30094b90300c289449619e9be98b827b619d4d7e8ddc460362949e9daeca7116;
  assign mdsMatrix_6_3 = 254'h2ad34bcfe341c5685c018acf0b5a7c11d9649534ca1e6c65c7432b4b0e646874;
  assign mdsMatrix_6_4 = 253'h173346c563ec6dbe554f8b0221dbfc5da410af5cce0f15e4949f788f1c24cfde;
  assign mdsMatrix_6_5 = 254'h284b46d9e6433e109fa41b53ef70ce50a47c184a41bda636d92727ec0fa535f8;
  assign mdsMatrix_6_6 = 253'h1922d0b4f4579c3a0b5009958af4264ba42544599875dcf9f6776366371a3321;
  assign mdsMatrix_6_7 = 254'h21a26b7357d55d3642edc6e9e7dacb31257897a5b5061594576285c95d709bda;
  assign mdsMatrix_6_8 = 254'h3dff06fa951718204dc2ba68d9ac05691d2e6652b1d2cb081395a535fc26aff8;
  assign mdsMatrix_6_9 = 254'h28e96e7538d3814f7ea7c94474969bb9b01017777f74aac9762028819aeb369f;
  assign mdsMatrix_6_10 = 255'h71b43412aa1ae069d402dbc23f8af7573d26601dbb047dd4d64b80e12a49514c;
  assign mdsMatrix_6_11 = 255'h40c549e33eea1bd9b1cc5fb2070f8c86f576e04cdfeda0c91698e118d32d3463;
  assign mdsMatrix_7_0 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_7_1 = 255'h5926065232ef9bedc453194039fc15e36da21887af005004ee3fd2cc28aef675;
  assign mdsMatrix_7_2 = 255'h41ee23f17d0025d61cd2578b9b47d8e2034c1999863c94b2b086e23a0c695685;
  assign mdsMatrix_7_3 = 255'h69d9f9f632557ac2c4ce207d2a80dc053bd63a7d505b1a8f93281484f38af5ba;
  assign mdsMatrix_7_4 = 254'h251e29d5bcec361c6a65da991cfb90f96f9f7c650bd94876f09fe8c9ab2c354c;
  assign mdsMatrix_7_5 = 253'h15064f004897e03209e30a2f225c50005d634ee8086ab971be720ed7339b8180;
  assign mdsMatrix_7_6 = 254'h21a26b7357d55d3642edc6e9e7dacb31257897a5b5061594576285c95d709bda;
  assign mdsMatrix_7_7 = 254'h3cc4bf5d76b740edf261f6ef772b48486e837c55bfed9be3087181f4540bb1de;
  assign mdsMatrix_7_8 = 253'h1ab79d87d85b0951eb9bc442e00f0ae80acd9b273b208ceaa09fca70a4ece8aa;
  assign mdsMatrix_7_9 = 255'h577c15fcbfa6feeb4f12823092efe2845b92c485660bbf17fbe2f055b58d90f8;
  assign mdsMatrix_7_10 = 255'h6dff1757db2872c5fdfd8cac63f186319ae62643c7730d65a559acdecc1f4641;
  assign mdsMatrix_7_11 = 255'h51dba391f014ee6462bbd49ad829dad346372ed2429c28e7760ca266764eaf64;
  assign mdsMatrix_8_0 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_8_1 = 255'h72a1062b57f4fa2e5771859d22f5fcd86130db83e0d506225b103cc5d3074aa7;
  assign mdsMatrix_8_2 = 254'h3cc52207bbd8577c030f4eb9521656c95a079c6c229005a7d5641c2e65c04144;
  assign mdsMatrix_8_3 = 255'h4177ffe5b5c4a55c525b37d5ec1f55eda6fade24205b20ba52cba1d4eb3d52b9;
  assign mdsMatrix_8_4 = 255'h4ebf8c6b40211b8a277d5a9d9d1014c18582596cf8ac3812e752af8428ba98e0;
  assign mdsMatrix_8_5 = 253'h1ae7d0b1501894960d8ef684c43bb9392c60c9f7c465d26081631de66ab866ef;
  assign mdsMatrix_8_6 = 254'h3dff06fa951718204dc2ba68d9ac05691d2e6652b1d2cb081395a535fc26aff8;
  assign mdsMatrix_8_7 = 253'h1ab79d87d85b0951eb9bc442e00f0ae80acd9b273b208ceaa09fca70a4ece8aa;
  assign mdsMatrix_8_8 = 255'h4fa374764d47eef86b98bcc83af630e76924dbc7be6850e3e52de26b1d5750bc;
  assign mdsMatrix_8_9 = 255'h68fc87287972d3ff6761576a7c69e0dc4eda93c9c53964688a1164e26d1ef4cf;
  assign mdsMatrix_8_10 = 255'h584b9a86f54718cf85eb1750395add2d56cde98fbfcb1aaa88224e105d0cd270;
  assign mdsMatrix_8_11 = 254'h3f7cd7bfb5918c72cc701a4a11d7271b76f46caed7a7f8823504df26f32aea61;
  assign mdsMatrix_9_0 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_9_1 = 254'h31d6995c6cfbe12818215b4349112482433988d1570f2c621c9e671a7684a3ef;
  assign mdsMatrix_9_2 = 254'h29ff2b59e1bc0353ecaf1d87cc085f91c8ed9b6212448aa1b5ceec55c996d003;
  assign mdsMatrix_9_3 = 255'h67e14645d098f70fa8c0e28a73bd0f75eceb766df2373013b1781684b482c9fb;
  assign mdsMatrix_9_4 = 254'h3ccfb0b82d30e2a96b4c21ed0cffffc34673eda2395e1b8db9cde8ab0e59d519;
  assign mdsMatrix_9_5 = 255'h4f6b915cd211c03922929e2bcda92d5d62c827224dbb0ec3ca13da4488dad173;
  assign mdsMatrix_9_6 = 254'h28e96e7538d3814f7ea7c94474969bb9b01017777f74aac9762028819aeb369f;
  assign mdsMatrix_9_7 = 255'h577c15fcbfa6feeb4f12823092efe2845b92c485660bbf17fbe2f055b58d90f8;
  assign mdsMatrix_9_8 = 255'h68fc87287972d3ff6761576a7c69e0dc4eda93c9c53964688a1164e26d1ef4cf;
  assign mdsMatrix_9_9 = 255'h62ada0082673eb09881466abf1fed60d2decf005ce699dc0f9963a0053a4f991;
  assign mdsMatrix_9_10 = 253'h15ba23b9eb93e2ea01b9e5f4bda6724acad35c979fd01d9e939b4d2a2e2a779a;
  assign mdsMatrix_9_11 = 254'h25ead4b041d15a5a823d731842893d31c82418c3d1ae98639b6059a78e11ad26;
  assign mdsMatrix_10_0 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_10_1 = 253'h14ff39ce71663ed6904498dc2b0cd2ffdd9f3da50d3b747d587adbd1ff4e192d;
  assign mdsMatrix_10_2 = 255'h5270a6310562c5907877e43b1bfa6e064ffdc02a8ec763fcf472d48e39acbd42;
  assign mdsMatrix_10_3 = 253'h197ba23e784e407b5d5513b59adbb98fa16dcb92bb6943197d3760b49b1dd1d1;
  assign mdsMatrix_10_4 = 253'h1ee8136953d9562ca3d0eb11698492c3c038b41c27d30886b5f4111f8a4e6c68;
  assign mdsMatrix_10_5 = 254'h2f9e31da3bca17f740ab3b2e13254875e6337da40fd7e6b76bfc9d776809c972;
  assign mdsMatrix_10_6 = 255'h71b43412aa1ae069d402dbc23f8af7573d26601dbb047dd4d64b80e12a49514c;
  assign mdsMatrix_10_7 = 255'h6dff1757db2872c5fdfd8cac63f186319ae62643c7730d65a559acdecc1f4641;
  assign mdsMatrix_10_8 = 255'h584b9a86f54718cf85eb1750395add2d56cde98fbfcb1aaa88224e105d0cd270;
  assign mdsMatrix_10_9 = 253'h15ba23b9eb93e2ea01b9e5f4bda6724acad35c979fd01d9e939b4d2a2e2a779a;
  assign mdsMatrix_10_10 = 255'h6d121e224aa9f67e2b13cd52bb37df74ed9e8aaaf7ef998efe0f7ecd3a1cb5a2;
  assign mdsMatrix_10_11 = 255'h501d48296076413d72abe7e778a8a98da6e6c7eeb020f3277b6f4fd7d1302058;
  assign mdsMatrix_11_0 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_11_1 = 255'h6a758500fad34882feffcb009873e6077e78d4300020f33ef22f40faba7981f7;
  assign mdsMatrix_11_2 = 254'h349cdd4bc00a305e5677872bbed238d65beae70b5f35522b3642560b63a5d7f0;
  assign mdsMatrix_11_3 = 255'h5753b589f9a06db49d750abe1351345af62a29ee5b6714168fc9785e6be004d3;
  assign mdsMatrix_11_4 = 255'h73a64e645c8c1cd18133f48ab3afdb4d1fae4241e83c6a4d429aa513f9a3414b;
  assign mdsMatrix_11_5 = 254'h39480b0425cd85cec7d8f43d000238cc3ca6805ba6fe7d8248330dc9bcdd1f18;
  assign mdsMatrix_11_6 = 255'h40c549e33eea1bd9b1cc5fb2070f8c86f576e04cdfeda0c91698e118d32d3463;
  assign mdsMatrix_11_7 = 255'h51dba391f014ee6462bbd49ad829dad346372ed2429c28e7760ca266764eaf64;
  assign mdsMatrix_11_8 = 254'h3f7cd7bfb5918c72cc701a4a11d7271b76f46caed7a7f8823504df26f32aea61;
  assign mdsMatrix_11_9 = 254'h25ead4b041d15a5a823d731842893d31c82418c3d1ae98639b6059a78e11ad26;
  assign mdsMatrix_11_10 = 255'h501d48296076413d72abe7e778a8a98da6e6c7eeb020f3277b6f4fd7d1302058;
  assign mdsMatrix_11_11 = 255'h664befc7faf5e8bf064497c2bdcff2241f3ccb9777045b67cd1353bdd8c345ac;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign tempAddrVec_5 = io_addr_regNext_5;
  assign tempAddrVec_6 = io_addr_regNext_6;
  assign tempAddrVec_7 = io_addr_regNext_7;
  assign tempAddrVec_8 = io_addr_regNext_8;
  assign tempAddrVec_9 = io_addr_regNext_9;
  assign tempAddrVec_10 = io_addr_regNext_10;
  assign tempAddrVec_11 = io_addr_regNext_11;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  assign io_data_5 = _zz_mdsMem_5_port0;
  assign io_data_6 = _zz_mdsMem_6_port0;
  assign io_data_7 = _zz_mdsMem_7_port0;
  assign io_data_8 = _zz_mdsMem_8_port0;
  assign io_data_9 = _zz_mdsMem_9_port0;
  assign io_data_10 = _zz_mdsMem_10_port0;
  assign io_data_11 = _zz_mdsMem_11_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
    io_addr_regNext_5 <= io_addr;
    io_addr_regNext_6 <= io_addr;
    io_addr_regNext_7 <= io_addr;
    io_addr_regNext_8 <= io_addr;
    io_addr_regNext_9 <= io_addr;
    io_addr_regNext_10 <= io_addr;
    io_addr_regNext_11 <= io_addr;
  end


endmodule

module MatrixConstantMem_6 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  input      [3:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  reg        [254:0]  _zz_mdsMem_5_port0;
  reg        [254:0]  _zz_mdsMem_6_port0;
  reg        [254:0]  _zz_mdsMem_7_port0;
  reg        [254:0]  _zz_mdsMem_8_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire                _zz_mdsMem_5_port;
  wire                _zz_io_data_5;
  wire                _zz_mdsMem_6_port;
  wire                _zz_io_data_6;
  wire                _zz_mdsMem_7_port;
  wire                _zz_io_data_7;
  wire                _zz_mdsMem_8_port;
  wire                _zz_io_data_8;
  wire       [254:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [253:0]  mdsMatrix_0_2;
  wire       [252:0]  mdsMatrix_0_3;
  wire       [254:0]  mdsMatrix_0_4;
  wire       [254:0]  mdsMatrix_0_5;
  wire       [252:0]  mdsMatrix_0_6;
  wire       [254:0]  mdsMatrix_0_7;
  wire       [253:0]  mdsMatrix_0_8;
  wire       [249:0]  mdsMatrix_1_0;
  wire       [247:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [254:0]  mdsMatrix_1_3;
  wire       [253:0]  mdsMatrix_1_4;
  wire       [254:0]  mdsMatrix_1_5;
  wire       [254:0]  mdsMatrix_1_6;
  wire       [253:0]  mdsMatrix_1_7;
  wire       [254:0]  mdsMatrix_1_8;
  wire       [253:0]  mdsMatrix_2_0;
  wire       [254:0]  mdsMatrix_2_1;
  wire       [254:0]  mdsMatrix_2_2;
  wire       [254:0]  mdsMatrix_2_3;
  wire       [254:0]  mdsMatrix_2_4;
  wire       [252:0]  mdsMatrix_2_5;
  wire       [254:0]  mdsMatrix_2_6;
  wire       [253:0]  mdsMatrix_2_7;
  wire       [254:0]  mdsMatrix_2_8;
  wire       [254:0]  mdsMatrix_3_0;
  wire       [254:0]  mdsMatrix_3_1;
  wire       [254:0]  mdsMatrix_3_2;
  wire       [253:0]  mdsMatrix_3_3;
  wire       [254:0]  mdsMatrix_3_4;
  wire       [254:0]  mdsMatrix_3_5;
  wire       [254:0]  mdsMatrix_3_6;
  wire       [253:0]  mdsMatrix_3_7;
  wire       [253:0]  mdsMatrix_3_8;
  wire       [254:0]  mdsMatrix_4_0;
  wire       [253:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [254:0]  mdsMatrix_4_3;
  wire       [253:0]  mdsMatrix_4_4;
  wire       [253:0]  mdsMatrix_4_5;
  wire       [254:0]  mdsMatrix_4_6;
  wire       [254:0]  mdsMatrix_4_7;
  wire       [254:0]  mdsMatrix_4_8;
  wire       [253:0]  mdsMatrix_5_0;
  wire       [254:0]  mdsMatrix_5_1;
  wire       [252:0]  mdsMatrix_5_2;
  wire       [254:0]  mdsMatrix_5_3;
  wire       [253:0]  mdsMatrix_5_4;
  wire       [253:0]  mdsMatrix_5_5;
  wire       [254:0]  mdsMatrix_5_6;
  wire       [253:0]  mdsMatrix_5_7;
  wire       [253:0]  mdsMatrix_5_8;
  wire       [254:0]  mdsMatrix_6_0;
  wire       [254:0]  mdsMatrix_6_1;
  wire       [254:0]  mdsMatrix_6_2;
  wire       [254:0]  mdsMatrix_6_3;
  wire       [254:0]  mdsMatrix_6_4;
  wire       [254:0]  mdsMatrix_6_5;
  wire       [253:0]  mdsMatrix_6_6;
  wire       [254:0]  mdsMatrix_6_7;
  wire       [253:0]  mdsMatrix_6_8;
  wire       [252:0]  mdsMatrix_7_0;
  wire       [253:0]  mdsMatrix_7_1;
  wire       [253:0]  mdsMatrix_7_2;
  wire       [253:0]  mdsMatrix_7_3;
  wire       [254:0]  mdsMatrix_7_4;
  wire       [253:0]  mdsMatrix_7_5;
  wire       [254:0]  mdsMatrix_7_6;
  wire       [254:0]  mdsMatrix_7_7;
  wire       [253:0]  mdsMatrix_7_8;
  wire       [253:0]  mdsMatrix_8_0;
  wire       [254:0]  mdsMatrix_8_1;
  wire       [254:0]  mdsMatrix_8_2;
  wire       [253:0]  mdsMatrix_8_3;
  wire       [254:0]  mdsMatrix_8_4;
  wire       [253:0]  mdsMatrix_8_5;
  wire       [253:0]  mdsMatrix_8_6;
  wire       [253:0]  mdsMatrix_8_7;
  wire       [253:0]  mdsMatrix_8_8;
  wire       [3:0]    tempAddrVec_0;
  wire       [3:0]    tempAddrVec_1;
  wire       [3:0]    tempAddrVec_2;
  wire       [3:0]    tempAddrVec_3;
  wire       [3:0]    tempAddrVec_4;
  wire       [3:0]    tempAddrVec_5;
  wire       [3:0]    tempAddrVec_6;
  wire       [3:0]    tempAddrVec_7;
  wire       [3:0]    tempAddrVec_8;
  reg        [3:0]    io_addr_regNext;
  reg        [3:0]    io_addr_regNext_1;
  reg        [3:0]    io_addr_regNext_2;
  reg        [3:0]    io_addr_regNext_3;
  reg        [3:0]    io_addr_regNext_4;
  reg        [3:0]    io_addr_regNext_5;
  reg        [3:0]    io_addr_regNext_6;
  reg        [3:0]    io_addr_regNext_7;
  reg        [3:0]    io_addr_regNext_8;
  reg [254:0] mdsMem_0 [0:8];
  reg [254:0] mdsMem_1 [0:8];
  reg [254:0] mdsMem_2 [0:8];
  reg [254:0] mdsMem_3 [0:8];
  reg [254:0] mdsMem_4 [0:8];
  reg [254:0] mdsMem_5 [0:8];
  reg [254:0] mdsMem_6 [0:8];
  reg [254:0] mdsMem_7 [0:8];
  reg [254:0] mdsMem_8 [0:8];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  assign _zz_io_data_5 = 1'b1;
  assign _zz_io_data_6 = 1'b1;
  assign _zz_io_data_7 = 1'b1;
  assign _zz_io_data_8 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_20_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_20_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_20_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_20_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_20_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_20_mdsMem_5.bin",mdsMem_5);
  end
  always @(posedge clk) begin
    if(_zz_io_data_5) begin
      _zz_mdsMem_5_port0 <= mdsMem_5[tempAddrVec_5];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_20_mdsMem_6.bin",mdsMem_6);
  end
  always @(posedge clk) begin
    if(_zz_io_data_6) begin
      _zz_mdsMem_6_port0 <= mdsMem_6[tempAddrVec_6];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_20_mdsMem_7.bin",mdsMem_7);
  end
  always @(posedge clk) begin
    if(_zz_io_data_7) begin
      _zz_mdsMem_7_port0 <= mdsMem_7[tempAddrVec_7];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_20_mdsMem_8.bin",mdsMem_8);
  end
  always @(posedge clk) begin
    if(_zz_io_data_8) begin
      _zz_mdsMem_8_port0 <= mdsMem_8[tempAddrVec_8];
    end
  end

  assign mdsMatrix_0_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_0_1 = 255'h5af7310f714af42f8111b0e51ccdecca129f01a21285bf4c0cf9b5092a09fadc;
  assign mdsMatrix_0_2 = 254'h2fcd74e4d241c2b43473b32b6d2b38713447261d83bec97c032c5dbcf589b4dc;
  assign mdsMatrix_0_3 = 253'h1377447987b7b82747f59b52e801efc237d95c4235013276442f4218edb98b25;
  assign mdsMatrix_0_4 = 255'h6ed258c11dd3e92f38525ad1e537213cc851dbe89595bf269415edce6f01ed3e;
  assign mdsMatrix_0_5 = 255'h6f32f1479a578cc93ed9cf1913cb21d5183aeafd6f47febde74a5597d8c01b72;
  assign mdsMatrix_0_6 = 253'h1330c90fbf4c108a82a9557731aacb7f5e0a46cded0f8eca84467ab8f8fede24;
  assign mdsMatrix_0_7 = 255'h5ec1004ffeeb5b19a368e25ceeb5d588ed7461e55a3afedf71e79cc72a958c54;
  assign mdsMatrix_0_8 = 254'h300a8b11d8240ad5a127153837de64677cb6ba792501065692fcbac4086dd7bc;
  assign mdsMatrix_1_0 = 250'h26a11bc2ae0808b28f46e64cadfa19888da1265cccd20cd0000000033333333;
  assign mdsMatrix_1_1 = 248'hc9e4b2f2574895016314e8e51e4dc0be2ce83ca40ba46fe9f48ec09eca2cbf;
  assign mdsMatrix_1_2 = 255'h6ca356aba3c6d3051810e5675865f34d344091d7e5f7130d1448e2da7c088254;
  assign mdsMatrix_1_3 = 255'h6bddeed58ed330235de0f187d5cd9ff4f55d249b8c68bad0111b052d2595f9cf;
  assign mdsMatrix_1_4 = 254'h38dcb36cb689adbfceab6bd2c66db3a312ac5c76920dfacf6489b8a6e57abf0d;
  assign mdsMatrix_1_5 = 255'h560c6b7a2173171bea8e4b372b9708591baf0793401516d6de46f093693e017d;
  assign mdsMatrix_1_6 = 255'h460fabe95f08dc6f86155fa415c298be3902451e7851890329f0e824951e4a40;
  assign mdsMatrix_1_7 = 254'h2329be65a7f8d6840673d3eef76939b4d69c99813404ba4588cac586ff1874f2;
  assign mdsMatrix_1_8 = 255'h62dcf8a2a99b248cf9eb57ece491381ca98d5a0f8bfaeef4544d0aa63d57a813;
  assign mdsMatrix_2_0 = 254'h2c59c154f04b2e0d209627474791ca2f8396d8008ba29c5ce8ba2e8b745d1746;
  assign mdsMatrix_2_1 = 255'h6ca356aba3c6d3051810e5675865f34d344091d7e5f7130d1448e2da7c088254;
  assign mdsMatrix_2_2 = 255'h4d8562d6924c0c936ba4ba7bf95520672783739c78cf1889302e81f3ce88277d;
  assign mdsMatrix_2_3 = 255'h6a5e9315e047b48bc8ad553d093fe5c4d07b15b468949f9ef169d01a7ab4ae15;
  assign mdsMatrix_2_4 = 255'h61c325e7484a00d30881b9495b7566790b14c9a85d2fb9499743cff01906e9f0;
  assign mdsMatrix_2_5 = 253'h13d974b3478565de14e3c8fb872bee0aed3b0aa662806d6d04bfe109db0365a0;
  assign mdsMatrix_2_6 = 255'h4aa47b9b992774232f36d89c24bb29bdf1a99654fc880181281dba2c3c4deba1;
  assign mdsMatrix_2_7 = 254'h2fae6443cfd4019977789b19c6041d7cada6d1b9683421b8e0ed05650ca875e5;
  assign mdsMatrix_2_8 = 255'h417490236aa5398ccabd839a416f1bd0895476ac32e8265fb2f8663445f55cba;
  assign mdsMatrix_3_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_3_1 = 255'h6bddeed58ed330235de0f187d5cd9ff4f55d249b8c68bad0111b052d2595f9cf;
  assign mdsMatrix_3_2 = 255'h6a5e9315e047b48bc8ad553d093fe5c4d07b15b468949f9ef169d01a7ab4ae15;
  assign mdsMatrix_3_3 = 254'h2c0bb77f030681e2867784a47cf698d97cbd73926dbf559d684fa66c48b6be4d;
  assign mdsMatrix_3_4 = 255'h56e0a9dff4e51ed01d2cbd39ab79a3ff2d800d0769807df87ae9d548a0b5c8db;
  assign mdsMatrix_3_5 = 255'h6d4b6fd9d7068dd8e3ce1a6b949e01a7f9ecbb6954d486c23ea79d928d31e1fb;
  assign mdsMatrix_3_6 = 255'h5d2f26a4e1e33d1353a7ae11a8312d4f7ba200af6bf977294df96acb19ff58ca;
  assign mdsMatrix_3_7 = 254'h289624559156d71b826b0f7df6aaf8e60e19845025682c0aba6d60b50022fdbd;
  assign mdsMatrix_3_8 = 254'h21653a9d03325193ffa49f4edd43af78fcbcd8677909e3147dc945c62762584f;
  assign mdsMatrix_4_0 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_4_1 = 254'h38dcb36cb689adbfceab6bd2c66db3a312ac5c76920dfacf6489b8a6e57abf0d;
  assign mdsMatrix_4_2 = 255'h61c325e7484a00d30881b9495b7566790b14c9a85d2fb9499743cff01906e9f0;
  assign mdsMatrix_4_3 = 255'h56e0a9dff4e51ed01d2cbd39ab79a3ff2d800d0769807df87ae9d548a0b5c8db;
  assign mdsMatrix_4_4 = 254'h3120e3b83a6f9e0c88e2210563d071ed564b3c2371f6ae12942da15cb4584fcc;
  assign mdsMatrix_4_5 = 254'h3d3fe7512e8c130a6183b760325dc21e6986c90556bcc099cda7ca87854186f5;
  assign mdsMatrix_4_6 = 255'h686e7728d8e7277f6871414c76d35956fbe54ed21cb5b6ba7843befddf7037c8;
  assign mdsMatrix_4_7 = 255'h4c63a6241edba92d3993229290be12b8a3ce8c593d10c3d6853f58fb207f58e3;
  assign mdsMatrix_4_8 = 255'h477c32cf4ff8ee74f62a432e68c0942216caff6c11bb17c081bb7f83856af896;
  assign mdsMatrix_5_0 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_5_1 = 255'h560c6b7a2173171bea8e4b372b9708591baf0793401516d6de46f093693e017d;
  assign mdsMatrix_5_2 = 253'h13d974b3478565de14e3c8fb872bee0aed3b0aa662806d6d04bfe109db0365a0;
  assign mdsMatrix_5_3 = 255'h6d4b6fd9d7068dd8e3ce1a6b949e01a7f9ecbb6954d486c23ea79d928d31e1fb;
  assign mdsMatrix_5_4 = 254'h3d3fe7512e8c130a6183b760325dc21e6986c90556bcc099cda7ca87854186f5;
  assign mdsMatrix_5_5 = 254'h2c271357a5bae475ea78679e98664012d84220ed2c5126fc6bd5770bf50915b1;
  assign mdsMatrix_5_6 = 255'h56f7569326d01da5966de3363569ea52a410477175bea44ef7b9d409e1c689c0;
  assign mdsMatrix_5_7 = 254'h3509f6a3a4ad7f83a9cca2e8c8232135d1d322f9233dff8cc089940843776d1c;
  assign mdsMatrix_5_8 = 254'h3cd8760ee40660f5934f465243213d0145de7d1874b7909f44e48785b2726dfa;
  assign mdsMatrix_6_0 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_6_1 = 255'h460fabe95f08dc6f86155fa415c298be3902451e7851890329f0e824951e4a40;
  assign mdsMatrix_6_2 = 255'h4aa47b9b992774232f36d89c24bb29bdf1a99654fc880181281dba2c3c4deba1;
  assign mdsMatrix_6_3 = 255'h5d2f26a4e1e33d1353a7ae11a8312d4f7ba200af6bf977294df96acb19ff58ca;
  assign mdsMatrix_6_4 = 255'h686e7728d8e7277f6871414c76d35956fbe54ed21cb5b6ba7843befddf7037c8;
  assign mdsMatrix_6_5 = 255'h56f7569326d01da5966de3363569ea52a410477175bea44ef7b9d409e1c689c0;
  assign mdsMatrix_6_6 = 254'h2897360218689ec9034dc0ca210c2c2e6cc480dd175d11f826f345abc8397257;
  assign mdsMatrix_6_7 = 255'h4cea8683dd9997312f53cc1d1e3dd066d2928df838c54e1c323fbbe605e484b6;
  assign mdsMatrix_6_8 = 254'h25424bca582695dad0cf15af89d6fff61cd3dedc995905886c2193acdad14ae7;
  assign mdsMatrix_7_0 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_7_1 = 254'h2329be65a7f8d6840673d3eef76939b4d69c99813404ba4588cac586ff1874f2;
  assign mdsMatrix_7_2 = 254'h2fae6443cfd4019977789b19c6041d7cada6d1b9683421b8e0ed05650ca875e5;
  assign mdsMatrix_7_3 = 254'h289624559156d71b826b0f7df6aaf8e60e19845025682c0aba6d60b50022fdbd;
  assign mdsMatrix_7_4 = 255'h4c63a6241edba92d3993229290be12b8a3ce8c593d10c3d6853f58fb207f58e3;
  assign mdsMatrix_7_5 = 254'h3509f6a3a4ad7f83a9cca2e8c8232135d1d322f9233dff8cc089940843776d1c;
  assign mdsMatrix_7_6 = 255'h4cea8683dd9997312f53cc1d1e3dd066d2928df838c54e1c323fbbe605e484b6;
  assign mdsMatrix_7_7 = 255'h5b0ea47c49e54a8949b5ac44bc4d03e7d6b3bdac7c5914a6cec40a74ae51a542;
  assign mdsMatrix_7_8 = 254'h3a5f57a8bf594bfc6e63cb3c9c4f4bea16c2790c3a678b58870ee149a5d1ac57;
  assign mdsMatrix_8_0 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_8_1 = 255'h62dcf8a2a99b248cf9eb57ece491381ca98d5a0f8bfaeef4544d0aa63d57a813;
  assign mdsMatrix_8_2 = 255'h417490236aa5398ccabd839a416f1bd0895476ac32e8265fb2f8663445f55cba;
  assign mdsMatrix_8_3 = 254'h21653a9d03325193ffa49f4edd43af78fcbcd8677909e3147dc945c62762584f;
  assign mdsMatrix_8_4 = 255'h477c32cf4ff8ee74f62a432e68c0942216caff6c11bb17c081bb7f83856af896;
  assign mdsMatrix_8_5 = 254'h3cd8760ee40660f5934f465243213d0145de7d1874b7909f44e48785b2726dfa;
  assign mdsMatrix_8_6 = 254'h25424bca582695dad0cf15af89d6fff61cd3dedc995905886c2193acdad14ae7;
  assign mdsMatrix_8_7 = 254'h3a5f57a8bf594bfc6e63cb3c9c4f4bea16c2790c3a678b58870ee149a5d1ac57;
  assign mdsMatrix_8_8 = 254'h36b3f71122dfee4322d02f20994fa1328e9146d146bf9569a2e945a460c82ee6;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign tempAddrVec_5 = io_addr_regNext_5;
  assign tempAddrVec_6 = io_addr_regNext_6;
  assign tempAddrVec_7 = io_addr_regNext_7;
  assign tempAddrVec_8 = io_addr_regNext_8;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  assign io_data_5 = _zz_mdsMem_5_port0;
  assign io_data_6 = _zz_mdsMem_6_port0;
  assign io_data_7 = _zz_mdsMem_7_port0;
  assign io_data_8 = _zz_mdsMem_8_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
    io_addr_regNext_5 <= io_addr;
    io_addr_regNext_6 <= io_addr;
    io_addr_regNext_7 <= io_addr;
    io_addr_regNext_8 <= io_addr;
  end


endmodule

module MatrixConstantMem_5 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  input      [2:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire       [250:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [253:0]  mdsMatrix_0_2;
  wire       [254:0]  mdsMatrix_0_3;
  wire       [254:0]  mdsMatrix_0_4;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [253:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [253:0]  mdsMatrix_1_3;
  wire       [252:0]  mdsMatrix_1_4;
  wire       [254:0]  mdsMatrix_2_0;
  wire       [254:0]  mdsMatrix_2_1;
  wire       [251:0]  mdsMatrix_2_2;
  wire       [252:0]  mdsMatrix_2_3;
  wire       [254:0]  mdsMatrix_2_4;
  wire       [253:0]  mdsMatrix_3_0;
  wire       [253:0]  mdsMatrix_3_1;
  wire       [252:0]  mdsMatrix_3_2;
  wire       [253:0]  mdsMatrix_3_3;
  wire       [252:0]  mdsMatrix_3_4;
  wire       [254:0]  mdsMatrix_4_0;
  wire       [252:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [252:0]  mdsMatrix_4_3;
  wire       [248:0]  mdsMatrix_4_4;
  wire       [2:0]    tempAddrVec_0;
  wire       [2:0]    tempAddrVec_1;
  wire       [2:0]    tempAddrVec_2;
  wire       [2:0]    tempAddrVec_3;
  wire       [2:0]    tempAddrVec_4;
  reg        [2:0]    io_addr_regNext;
  reg        [2:0]    io_addr_regNext_1;
  reg        [2:0]    io_addr_regNext_2;
  reg        [2:0]    io_addr_regNext_3;
  reg        [2:0]    io_addr_regNext_4;
  reg [254:0] mdsMem_0 [0:4];
  reg [254:0] mdsMem_1 [0:4];
  reg [254:0] mdsMem_2 [0:4];
  reg [254:0] mdsMem_3 [0:4];
  reg [254:0] mdsMem_4 [0:4];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_19_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_19_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_19_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_19_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_19_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  assign mdsMatrix_0_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_0_1 = 255'h5301f64426b3ebca1f6651d78d256903f80141c43c2e8f2d5c42429d2da832c9;
  assign mdsMatrix_0_2 = 254'h3d7e2fe8a9cf4c482ad7e335060ee024ab7c02cdee8d79c488bc776a7277500d;
  assign mdsMatrix_0_3 = 255'h5fb37b8083eeb410ed792f28064ab12da369d8c6ea8f3b11bdf953ecf125f70c;
  assign mdsMatrix_0_4 = 255'h57fabbc58de3cee7b6c5f61d7399f980b41ff9e0c1fc4099ae0f225c901e444d;
  assign mdsMatrix_1_0 = 255'h514f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_1_1 = 254'h3b13122516ea9c45f99cec6182cd8f49d4ecba0ec0fa58c132342950ee316a69;
  assign mdsMatrix_1_2 = 255'h48b3669cc94450051fbb37f9a37576dcf43f7419c9e80d8d1b55c267d36851b4;
  assign mdsMatrix_1_3 = 254'h29386bc84ccab5b73cd7f602762aed1b2db36d3d0ef1f77134c8e7f44874c4d3;
  assign mdsMatrix_1_4 = 253'h1b1a2fb021ae315d87c4202ad51ea54ed8429784720de9ac59ed11f884f9c9c7;
  assign mdsMatrix_2_0 = 255'h66d0f1e660ec4796f8b356e005810db9e6b5824adb6cc6dadb6db6dadb6db6dc;
  assign mdsMatrix_2_1 = 255'h48b3669cc94450051fbb37f9a37576dcf43f7419c9e80d8d1b55c267d36851b4;
  assign mdsMatrix_2_2 = 252'hc3f3140031a893bbfdc443c2786c6518ca6690d226ef7d333d42512ff3720cc;
  assign mdsMatrix_2_3 = 253'h1f0c1edd5e10ea8b940df709c813ff880e4fac115efe0113554907b997612380;
  assign mdsMatrix_2_4 = 255'h5e35a96c7dfa83af31d6ea2882e74655589a02c86410f5b0e58fd0c8599858a6;
  assign mdsMatrix_3_0 = 254'h2000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_3_1 = 254'h29386bc84ccab5b73cd7f602762aed1b2db36d3d0ef1f77134c8e7f44874c4d3;
  assign mdsMatrix_3_2 = 253'h1f0c1edd5e10ea8b940df709c813ff880e4fac115efe0113554907b997612380;
  assign mdsMatrix_3_3 = 254'h2e3e6a432b5b0226ce6f0e65b1d20e5434b4072d7e4733208d7b739051aab926;
  assign mdsMatrix_3_4 = 253'h14769e2082dd9a34a211d4fe8e8e097a66d1c33bd4e22affbb6133ddfc5fcf30;
  assign mdsMatrix_4_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_4_1 = 253'h1b1a2fb021ae315d87c4202ad51ea54ed8429784720de9ac59ed11f884f9c9c7;
  assign mdsMatrix_4_2 = 255'h5e35a96c7dfa83af31d6ea2882e74655589a02c86410f5b0e58fd0c8599858a6;
  assign mdsMatrix_4_3 = 253'h14769e2082dd9a34a211d4fe8e8e097a66d1c33bd4e22affbb6133ddfc5fcf30;
  assign mdsMatrix_4_4 = 249'h1d11e38f8014a70be5c6e4c025773b9ef6649d8ceb30ddb2492c459085fc174;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
  end


endmodule

module MatrixConstantMem_4 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  input      [1:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire       [253:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [253:0]  mdsMatrix_0_2;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [254:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [250:0]  mdsMatrix_2_0;
  wire       [254:0]  mdsMatrix_2_1;
  wire       [252:0]  mdsMatrix_2_2;
  wire       [1:0]    tempAddrVec_0;
  wire       [1:0]    tempAddrVec_1;
  wire       [1:0]    tempAddrVec_2;
  reg        [1:0]    io_addr_regNext;
  reg        [1:0]    io_addr_regNext_1;
  reg        [1:0]    io_addr_regNext_2;
  reg [254:0] mdsMem_0 [0:2];
  reg [254:0] mdsMem_1 [0:2];
  reg [254:0] mdsMem_2 [0:2];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_18_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_18_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_18_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  assign mdsMatrix_0_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_0_1 = 255'h516cfbe5a0499eb26e0db7e149cb1614f2159006be9dd597e7ad644f2cc8fcce;
  assign mdsMatrix_0_2 = 254'h2b5d8fedce156062b41e31b3e4051fb39def47675840ccfd40b77fb2a5c1dcc6;
  assign mdsMatrix_1_0 = 255'h4000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_1_1 = 255'h717f183d735a42a911080d993a296f1bdc192f9a7c8a38d8a4e176e6b856e237;
  assign mdsMatrix_1_2 = 255'h65483579139538bf910625005ee03a4d92a041b4572547b064d724c2907def5a;
  assign mdsMatrix_2_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_2_1 = 255'h65483579139538bf910625005ee03a4d92a041b4572547b064d724c2907def5a;
  assign mdsMatrix_2_2 = 253'h1326a139a061135832adaf114f318cefe528f09cf0f3500a650cbac1c8a0bc09;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
  end


endmodule

module MatrixConstantMem_3 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  output     [254:0]  io_data_9,
  output     [254:0]  io_data_10,
  output     [254:0]  io_data_11,
  input      [3:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  reg        [254:0]  _zz_mdsMem_5_port0;
  reg        [254:0]  _zz_mdsMem_6_port0;
  reg        [254:0]  _zz_mdsMem_7_port0;
  reg        [254:0]  _zz_mdsMem_8_port0;
  reg        [254:0]  _zz_mdsMem_9_port0;
  reg        [254:0]  _zz_mdsMem_10_port0;
  reg        [254:0]  _zz_mdsMem_11_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire                _zz_mdsMem_5_port;
  wire                _zz_io_data_5;
  wire                _zz_mdsMem_6_port;
  wire                _zz_io_data_6;
  wire                _zz_mdsMem_7_port;
  wire                _zz_io_data_7;
  wire                _zz_mdsMem_8_port;
  wire                _zz_io_data_8;
  wire                _zz_mdsMem_9_port;
  wire                _zz_io_data_9;
  wire                _zz_mdsMem_10_port;
  wire                _zz_io_data_10;
  wire                _zz_mdsMem_11_port;
  wire                _zz_io_data_11;
  wire       [254:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [253:0]  mdsMatrix_0_2;
  wire       [254:0]  mdsMatrix_0_3;
  wire       [252:0]  mdsMatrix_0_4;
  wire       [253:0]  mdsMatrix_0_5;
  wire       [254:0]  mdsMatrix_0_6;
  wire       [252:0]  mdsMatrix_0_7;
  wire       [253:0]  mdsMatrix_0_8;
  wire       [254:0]  mdsMatrix_0_9;
  wire       [252:0]  mdsMatrix_0_10;
  wire       [250:0]  mdsMatrix_0_11;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [253:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [252:0]  mdsMatrix_1_3;
  wire       [253:0]  mdsMatrix_1_4;
  wire       [254:0]  mdsMatrix_1_5;
  wire       [252:0]  mdsMatrix_1_6;
  wire       [253:0]  mdsMatrix_1_7;
  wire       [254:0]  mdsMatrix_1_8;
  wire       [252:0]  mdsMatrix_1_9;
  wire       [250:0]  mdsMatrix_1_10;
  wire       [253:0]  mdsMatrix_1_11;
  wire       [253:0]  mdsMatrix_2_0;
  wire       [254:0]  mdsMatrix_2_1;
  wire       [252:0]  mdsMatrix_2_2;
  wire       [253:0]  mdsMatrix_2_3;
  wire       [254:0]  mdsMatrix_2_4;
  wire       [252:0]  mdsMatrix_2_5;
  wire       [253:0]  mdsMatrix_2_6;
  wire       [254:0]  mdsMatrix_2_7;
  wire       [252:0]  mdsMatrix_2_8;
  wire       [250:0]  mdsMatrix_2_9;
  wire       [253:0]  mdsMatrix_2_10;
  wire       [252:0]  mdsMatrix_2_11;
  wire       [254:0]  mdsMatrix_3_0;
  wire       [252:0]  mdsMatrix_3_1;
  wire       [253:0]  mdsMatrix_3_2;
  wire       [254:0]  mdsMatrix_3_3;
  wire       [252:0]  mdsMatrix_3_4;
  wire       [253:0]  mdsMatrix_3_5;
  wire       [254:0]  mdsMatrix_3_6;
  wire       [252:0]  mdsMatrix_3_7;
  wire       [250:0]  mdsMatrix_3_8;
  wire       [253:0]  mdsMatrix_3_9;
  wire       [252:0]  mdsMatrix_3_10;
  wire       [254:0]  mdsMatrix_3_11;
  wire       [252:0]  mdsMatrix_4_0;
  wire       [253:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [252:0]  mdsMatrix_4_3;
  wire       [253:0]  mdsMatrix_4_4;
  wire       [254:0]  mdsMatrix_4_5;
  wire       [252:0]  mdsMatrix_4_6;
  wire       [250:0]  mdsMatrix_4_7;
  wire       [253:0]  mdsMatrix_4_8;
  wire       [252:0]  mdsMatrix_4_9;
  wire       [254:0]  mdsMatrix_4_10;
  wire       [252:0]  mdsMatrix_4_11;
  wire       [253:0]  mdsMatrix_5_0;
  wire       [254:0]  mdsMatrix_5_1;
  wire       [252:0]  mdsMatrix_5_2;
  wire       [253:0]  mdsMatrix_5_3;
  wire       [254:0]  mdsMatrix_5_4;
  wire       [252:0]  mdsMatrix_5_5;
  wire       [250:0]  mdsMatrix_5_6;
  wire       [253:0]  mdsMatrix_5_7;
  wire       [252:0]  mdsMatrix_5_8;
  wire       [254:0]  mdsMatrix_5_9;
  wire       [252:0]  mdsMatrix_5_10;
  wire       [252:0]  mdsMatrix_5_11;
  wire       [254:0]  mdsMatrix_6_0;
  wire       [252:0]  mdsMatrix_6_1;
  wire       [253:0]  mdsMatrix_6_2;
  wire       [254:0]  mdsMatrix_6_3;
  wire       [252:0]  mdsMatrix_6_4;
  wire       [250:0]  mdsMatrix_6_5;
  wire       [253:0]  mdsMatrix_6_6;
  wire       [252:0]  mdsMatrix_6_7;
  wire       [254:0]  mdsMatrix_6_8;
  wire       [252:0]  mdsMatrix_6_9;
  wire       [252:0]  mdsMatrix_6_10;
  wire       [254:0]  mdsMatrix_6_11;
  wire       [252:0]  mdsMatrix_7_0;
  wire       [253:0]  mdsMatrix_7_1;
  wire       [254:0]  mdsMatrix_7_2;
  wire       [252:0]  mdsMatrix_7_3;
  wire       [250:0]  mdsMatrix_7_4;
  wire       [253:0]  mdsMatrix_7_5;
  wire       [252:0]  mdsMatrix_7_6;
  wire       [254:0]  mdsMatrix_7_7;
  wire       [252:0]  mdsMatrix_7_8;
  wire       [252:0]  mdsMatrix_7_9;
  wire       [254:0]  mdsMatrix_7_10;
  wire       [253:0]  mdsMatrix_7_11;
  wire       [253:0]  mdsMatrix_8_0;
  wire       [254:0]  mdsMatrix_8_1;
  wire       [252:0]  mdsMatrix_8_2;
  wire       [250:0]  mdsMatrix_8_3;
  wire       [253:0]  mdsMatrix_8_4;
  wire       [252:0]  mdsMatrix_8_5;
  wire       [254:0]  mdsMatrix_8_6;
  wire       [252:0]  mdsMatrix_8_7;
  wire       [252:0]  mdsMatrix_8_8;
  wire       [254:0]  mdsMatrix_8_9;
  wire       [253:0]  mdsMatrix_8_10;
  wire       [254:0]  mdsMatrix_8_11;
  wire       [254:0]  mdsMatrix_9_0;
  wire       [252:0]  mdsMatrix_9_1;
  wire       [250:0]  mdsMatrix_9_2;
  wire       [253:0]  mdsMatrix_9_3;
  wire       [252:0]  mdsMatrix_9_4;
  wire       [254:0]  mdsMatrix_9_5;
  wire       [252:0]  mdsMatrix_9_6;
  wire       [252:0]  mdsMatrix_9_7;
  wire       [254:0]  mdsMatrix_9_8;
  wire       [253:0]  mdsMatrix_9_9;
  wire       [254:0]  mdsMatrix_9_10;
  wire       [251:0]  mdsMatrix_9_11;
  wire       [252:0]  mdsMatrix_10_0;
  wire       [250:0]  mdsMatrix_10_1;
  wire       [253:0]  mdsMatrix_10_2;
  wire       [252:0]  mdsMatrix_10_3;
  wire       [254:0]  mdsMatrix_10_4;
  wire       [252:0]  mdsMatrix_10_5;
  wire       [252:0]  mdsMatrix_10_6;
  wire       [254:0]  mdsMatrix_10_7;
  wire       [253:0]  mdsMatrix_10_8;
  wire       [254:0]  mdsMatrix_10_9;
  wire       [251:0]  mdsMatrix_10_10;
  wire       [251:0]  mdsMatrix_10_11;
  wire       [250:0]  mdsMatrix_11_0;
  wire       [253:0]  mdsMatrix_11_1;
  wire       [252:0]  mdsMatrix_11_2;
  wire       [254:0]  mdsMatrix_11_3;
  wire       [252:0]  mdsMatrix_11_4;
  wire       [252:0]  mdsMatrix_11_5;
  wire       [254:0]  mdsMatrix_11_6;
  wire       [253:0]  mdsMatrix_11_7;
  wire       [254:0]  mdsMatrix_11_8;
  wire       [251:0]  mdsMatrix_11_9;
  wire       [251:0]  mdsMatrix_11_10;
  wire       [252:0]  mdsMatrix_11_11;
  wire       [3:0]    tempAddrVec_0;
  wire       [3:0]    tempAddrVec_1;
  wire       [3:0]    tempAddrVec_2;
  wire       [3:0]    tempAddrVec_3;
  wire       [3:0]    tempAddrVec_4;
  wire       [3:0]    tempAddrVec_5;
  wire       [3:0]    tempAddrVec_6;
  wire       [3:0]    tempAddrVec_7;
  wire       [3:0]    tempAddrVec_8;
  wire       [3:0]    tempAddrVec_9;
  wire       [3:0]    tempAddrVec_10;
  wire       [3:0]    tempAddrVec_11;
  reg        [3:0]    io_addr_regNext;
  reg        [3:0]    io_addr_regNext_1;
  reg        [3:0]    io_addr_regNext_2;
  reg        [3:0]    io_addr_regNext_3;
  reg        [3:0]    io_addr_regNext_4;
  reg        [3:0]    io_addr_regNext_5;
  reg        [3:0]    io_addr_regNext_6;
  reg        [3:0]    io_addr_regNext_7;
  reg        [3:0]    io_addr_regNext_8;
  reg        [3:0]    io_addr_regNext_9;
  reg        [3:0]    io_addr_regNext_10;
  reg        [3:0]    io_addr_regNext_11;
  reg [254:0] mdsMem_0 [0:11];
  reg [254:0] mdsMem_1 [0:11];
  reg [254:0] mdsMem_2 [0:11];
  reg [254:0] mdsMem_3 [0:11];
  reg [254:0] mdsMem_4 [0:11];
  reg [254:0] mdsMem_5 [0:11];
  reg [254:0] mdsMem_6 [0:11];
  reg [254:0] mdsMem_7 [0:11];
  reg [254:0] mdsMem_8 [0:11];
  reg [254:0] mdsMem_9 [0:11];
  reg [254:0] mdsMem_10 [0:11];
  reg [254:0] mdsMem_11 [0:11];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  assign _zz_io_data_5 = 1'b1;
  assign _zz_io_data_6 = 1'b1;
  assign _zz_io_data_7 = 1'b1;
  assign _zz_io_data_8 = 1'b1;
  assign _zz_io_data_9 = 1'b1;
  assign _zz_io_data_10 = 1'b1;
  assign _zz_io_data_11 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_5.bin",mdsMem_5);
  end
  always @(posedge clk) begin
    if(_zz_io_data_5) begin
      _zz_mdsMem_5_port0 <= mdsMem_5[tempAddrVec_5];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_6.bin",mdsMem_6);
  end
  always @(posedge clk) begin
    if(_zz_io_data_6) begin
      _zz_mdsMem_6_port0 <= mdsMem_6[tempAddrVec_6];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_7.bin",mdsMem_7);
  end
  always @(posedge clk) begin
    if(_zz_io_data_7) begin
      _zz_mdsMem_7_port0 <= mdsMem_7[tempAddrVec_7];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_8.bin",mdsMem_8);
  end
  always @(posedge clk) begin
    if(_zz_io_data_8) begin
      _zz_mdsMem_8_port0 <= mdsMem_8[tempAddrVec_8];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_9.bin",mdsMem_9);
  end
  always @(posedge clk) begin
    if(_zz_io_data_9) begin
      _zz_mdsMem_9_port0 <= mdsMem_9[tempAddrVec_9];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_10.bin",mdsMem_10);
  end
  always @(posedge clk) begin
    if(_zz_io_data_10) begin
      _zz_mdsMem_10_port0 <= mdsMem_10[tempAddrVec_10];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_17_mdsMem_11.bin",mdsMem_11);
  end
  always @(posedge clk) begin
    if(_zz_io_data_11) begin
      _zz_mdsMem_11_port0 <= mdsMem_11[tempAddrVec_11];
    end
  end

  assign mdsMatrix_0_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_0_1 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_0_2 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_0_3 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_0_4 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_0_5 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_0_6 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_0_7 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_0_8 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_0_9 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_0_10 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_0_11 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_1_0 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_1_1 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_1_2 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_1_3 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_1_4 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_1_5 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_1_6 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_1_7 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_1_8 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_1_9 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_1_10 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_1_11 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_2_0 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_2_1 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_2_2 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_2_3 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_2_4 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_2_5 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_2_6 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_2_7 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_2_8 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_2_9 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_2_10 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_2_11 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_3_0 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_3_1 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_3_2 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_3_3 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_3_4 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_3_5 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_3_6 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_3_7 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_3_8 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_3_9 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_3_10 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_3_11 = 255'h630594675b16af23d8a2a62d91416b17ca431bb389d75a7562762761b13b13b2;
  assign mdsMatrix_4_0 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_4_1 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_4_2 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_4_3 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_4_4 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_4_5 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_4_6 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_4_7 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_4_8 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_4_9 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_4_10 = 255'h630594675b16af23d8a2a62d91416b17ca431bb389d75a7562762761b13b13b2;
  assign mdsMatrix_4_11 = 253'h1ef31efc7000b862b42728017d0b0213f31027daa12f1a848e38e38e097b425f;
  assign mdsMatrix_5_0 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_5_1 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_5_2 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_5_3 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_5_4 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_5_5 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_5_6 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_5_7 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_5_8 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_5_9 = 255'h630594675b16af23d8a2a62d91416b17ca431bb389d75a7562762761b13b13b2;
  assign mdsMatrix_5_10 = 253'h1ef31efc7000b862b42728017d0b0213f31027daa12f1a848e38e38e097b425f;
  assign mdsMatrix_5_11 = 253'h19b43c79983b11e5be2cd5b80160436e79ad6092b6db31b6b6db6db6b6db6db7;
  assign mdsMatrix_6_0 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_6_1 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_6_2 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_6_3 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_6_4 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_6_5 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_6_6 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_6_7 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_6_8 = 255'h630594675b16af23d8a2a62d91416b17ca431bb389d75a7562762761b13b13b2;
  assign mdsMatrix_6_9 = 253'h1ef31efc7000b862b42728017d0b0213f31027daa12f1a848e38e38e097b425f;
  assign mdsMatrix_6_10 = 253'h19b43c79983b11e5be2cd5b80160436e79ad6092b6db31b6b6db6db6b6db6db7;
  assign mdsMatrix_6_11 = 255'h70c369e0a0e579263f94f6a61a4a7b0d9a86b65af72aaac14f72c23411a7b962;
  assign mdsMatrix_7_0 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_7_1 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_7_2 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_7_3 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_7_4 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_7_5 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_7_6 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_7_7 = 255'h630594675b16af23d8a2a62d91416b17ca431bb389d75a7562762761b13b13b2;
  assign mdsMatrix_7_8 = 253'h1ef31efc7000b862b42728017d0b0213f31027daa12f1a848e38e38e097b425f;
  assign mdsMatrix_7_9 = 253'h19b43c79983b11e5be2cd5b80160436e79ad6092b6db31b6b6db6db6b6db6db7;
  assign mdsMatrix_7_10 = 255'h70c369e0a0e579263f94f6a61a4a7b0d9a86b65af72aaac14f72c23411a7b962;
  assign mdsMatrix_7_11 = 254'h277293051c29ff46740f6ccef1807ddf4987e7784443d443ffffffffbbbbbbbc;
  assign mdsMatrix_8_0 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_8_1 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_8_2 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_8_3 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_8_4 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_8_5 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_8_6 = 255'h630594675b16af23d8a2a62d91416b17ca431bb389d75a7562762761b13b13b2;
  assign mdsMatrix_8_7 = 253'h1ef31efc7000b862b42728017d0b0213f31027daa12f1a848e38e38e097b425f;
  assign mdsMatrix_8_8 = 253'h19b43c79983b11e5be2cd5b80160436e79ad6092b6db31b6b6db6db6b6db6db7;
  assign mdsMatrix_8_9 = 255'h70c369e0a0e579263f94f6a61a4a7b0d9a86b65af72aaac14f72c23411a7b962;
  assign mdsMatrix_8_10 = 254'h277293051c29ff46740f6ccef1807ddf4987e7784443d443ffffffffbbbbbbbc;
  assign mdsMatrix_8_11 = 255'h4b92401fc595407c80d743a191fae08738e1ba12420f90417bdef7bd5ad6b5ae;
  assign mdsMatrix_9_0 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_9_1 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_9_2 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_9_3 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_9_4 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_9_5 = 255'h630594675b16af23d8a2a62d91416b17ca431bb389d75a7562762761b13b13b2;
  assign mdsMatrix_9_6 = 253'h1ef31efc7000b862b42728017d0b0213f31027daa12f1a848e38e38e097b425f;
  assign mdsMatrix_9_7 = 253'h19b43c79983b11e5be2cd5b80160436e79ad6092b6db31b6b6db6db6b6db6db7;
  assign mdsMatrix_9_8 = 255'h70c369e0a0e579263f94f6a61a4a7b0d9a86b65af72aaac14f72c23411a7b962;
  assign mdsMatrix_9_9 = 254'h277293051c29ff46740f6ccef1807ddf4987e7784443d443ffffffffbbbbbbbc;
  assign mdsMatrix_9_10 = 255'h4b92401fc595407c80d743a191fae08738e1ba12420f90417bdef7bd5ad6b5ae;
  assign mdsMatrix_9_11 = 252'h800000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_10_0 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_10_1 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_10_2 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_10_3 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_10_4 = 255'h630594675b16af23d8a2a62d91416b17ca431bb389d75a7562762761b13b13b2;
  assign mdsMatrix_10_5 = 253'h1ef31efc7000b862b42728017d0b0213f31027daa12f1a848e38e38e097b425f;
  assign mdsMatrix_10_6 = 253'h19b43c79983b11e5be2cd5b80160436e79ad6092b6db31b6b6db6db6b6db6db7;
  assign mdsMatrix_10_7 = 255'h70c369e0a0e579263f94f6a61a4a7b0d9a86b65af72aaac14f72c23411a7b962;
  assign mdsMatrix_10_8 = 254'h277293051c29ff46740f6ccef1807ddf4987e7784443d443ffffffffbbbbbbbc;
  assign mdsMatrix_10_9 = 255'h4b92401fc595407c80d743a191fae08738e1ba12420f90417bdef7bd5ad6b5ae;
  assign mdsMatrix_10_10 = 252'h800000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_10_11 = 252'hec895c6fac3ba0460320d17c285ee0fd6879d5583e0dec9a2e8ba2e7c1f07c2;
  assign mdsMatrix_11_0 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_11_1 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_11_2 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign mdsMatrix_11_3 = 255'h630594675b16af23d8a2a62d91416b17ca431bb389d75a7562762761b13b13b2;
  assign mdsMatrix_11_4 = 253'h1ef31efc7000b862b42728017d0b0213f31027daa12f1a848e38e38e097b425f;
  assign mdsMatrix_11_5 = 253'h19b43c79983b11e5be2cd5b80160436e79ad6092b6db31b6b6db6db6b6db6db7;
  assign mdsMatrix_11_6 = 255'h70c369e0a0e579263f94f6a61a4a7b0d9a86b65af72aaac14f72c23411a7b962;
  assign mdsMatrix_11_7 = 254'h277293051c29ff46740f6ccef1807ddf4987e7784443d443ffffffffbbbbbbbc;
  assign mdsMatrix_11_8 = 255'h4b92401fc595407c80d743a191fae08738e1ba12420f90417bdef7bd5ad6b5ae;
  assign mdsMatrix_11_9 = 252'h800000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_11_10 = 252'hec895c6fac3ba0460320d17c285ee0fd6879d5583e0dec9a2e8ba2e7c1f07c2;
  assign mdsMatrix_11_11 = 253'h152b04a05f3fb462d8d9a0f1e303fb4bebbbf52d8787561dffffffffe1e1e1e2;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign tempAddrVec_5 = io_addr_regNext_5;
  assign tempAddrVec_6 = io_addr_regNext_6;
  assign tempAddrVec_7 = io_addr_regNext_7;
  assign tempAddrVec_8 = io_addr_regNext_8;
  assign tempAddrVec_9 = io_addr_regNext_9;
  assign tempAddrVec_10 = io_addr_regNext_10;
  assign tempAddrVec_11 = io_addr_regNext_11;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  assign io_data_5 = _zz_mdsMem_5_port0;
  assign io_data_6 = _zz_mdsMem_6_port0;
  assign io_data_7 = _zz_mdsMem_7_port0;
  assign io_data_8 = _zz_mdsMem_8_port0;
  assign io_data_9 = _zz_mdsMem_9_port0;
  assign io_data_10 = _zz_mdsMem_10_port0;
  assign io_data_11 = _zz_mdsMem_11_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
    io_addr_regNext_5 <= io_addr;
    io_addr_regNext_6 <= io_addr;
    io_addr_regNext_7 <= io_addr;
    io_addr_regNext_8 <= io_addr;
    io_addr_regNext_9 <= io_addr;
    io_addr_regNext_10 <= io_addr;
    io_addr_regNext_11 <= io_addr;
  end


endmodule

module MatrixConstantMem_2 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  output     [254:0]  io_data_5,
  output     [254:0]  io_data_6,
  output     [254:0]  io_data_7,
  output     [254:0]  io_data_8,
  input      [3:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  reg        [254:0]  _zz_mdsMem_5_port0;
  reg        [254:0]  _zz_mdsMem_6_port0;
  reg        [254:0]  _zz_mdsMem_7_port0;
  reg        [254:0]  _zz_mdsMem_8_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire                _zz_mdsMem_5_port;
  wire                _zz_io_data_5;
  wire                _zz_mdsMem_6_port;
  wire                _zz_io_data_6;
  wire                _zz_mdsMem_7_port;
  wire                _zz_io_data_7;
  wire                _zz_mdsMem_8_port;
  wire                _zz_io_data_8;
  wire       [254:0]  mdsMatrix_0_0;
  wire       [249:0]  mdsMatrix_0_1;
  wire       [253:0]  mdsMatrix_0_2;
  wire       [254:0]  mdsMatrix_0_3;
  wire       [254:0]  mdsMatrix_0_4;
  wire       [253:0]  mdsMatrix_0_5;
  wire       [254:0]  mdsMatrix_0_6;
  wire       [252:0]  mdsMatrix_0_7;
  wire       [253:0]  mdsMatrix_0_8;
  wire       [249:0]  mdsMatrix_1_0;
  wire       [253:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [254:0]  mdsMatrix_1_3;
  wire       [253:0]  mdsMatrix_1_4;
  wire       [254:0]  mdsMatrix_1_5;
  wire       [252:0]  mdsMatrix_1_6;
  wire       [253:0]  mdsMatrix_1_7;
  wire       [254:0]  mdsMatrix_1_8;
  wire       [253:0]  mdsMatrix_2_0;
  wire       [254:0]  mdsMatrix_2_1;
  wire       [254:0]  mdsMatrix_2_2;
  wire       [253:0]  mdsMatrix_2_3;
  wire       [254:0]  mdsMatrix_2_4;
  wire       [252:0]  mdsMatrix_2_5;
  wire       [253:0]  mdsMatrix_2_6;
  wire       [254:0]  mdsMatrix_2_7;
  wire       [252:0]  mdsMatrix_2_8;
  wire       [254:0]  mdsMatrix_3_0;
  wire       [254:0]  mdsMatrix_3_1;
  wire       [253:0]  mdsMatrix_3_2;
  wire       [254:0]  mdsMatrix_3_3;
  wire       [252:0]  mdsMatrix_3_4;
  wire       [253:0]  mdsMatrix_3_5;
  wire       [254:0]  mdsMatrix_3_6;
  wire       [252:0]  mdsMatrix_3_7;
  wire       [253:0]  mdsMatrix_3_8;
  wire       [254:0]  mdsMatrix_4_0;
  wire       [253:0]  mdsMatrix_4_1;
  wire       [254:0]  mdsMatrix_4_2;
  wire       [252:0]  mdsMatrix_4_3;
  wire       [253:0]  mdsMatrix_4_4;
  wire       [254:0]  mdsMatrix_4_5;
  wire       [252:0]  mdsMatrix_4_6;
  wire       [253:0]  mdsMatrix_4_7;
  wire       [254:0]  mdsMatrix_4_8;
  wire       [253:0]  mdsMatrix_5_0;
  wire       [254:0]  mdsMatrix_5_1;
  wire       [252:0]  mdsMatrix_5_2;
  wire       [253:0]  mdsMatrix_5_3;
  wire       [254:0]  mdsMatrix_5_4;
  wire       [252:0]  mdsMatrix_5_5;
  wire       [253:0]  mdsMatrix_5_6;
  wire       [254:0]  mdsMatrix_5_7;
  wire       [252:0]  mdsMatrix_5_8;
  wire       [254:0]  mdsMatrix_6_0;
  wire       [252:0]  mdsMatrix_6_1;
  wire       [253:0]  mdsMatrix_6_2;
  wire       [254:0]  mdsMatrix_6_3;
  wire       [252:0]  mdsMatrix_6_4;
  wire       [253:0]  mdsMatrix_6_5;
  wire       [254:0]  mdsMatrix_6_6;
  wire       [252:0]  mdsMatrix_6_7;
  wire       [250:0]  mdsMatrix_6_8;
  wire       [252:0]  mdsMatrix_7_0;
  wire       [253:0]  mdsMatrix_7_1;
  wire       [254:0]  mdsMatrix_7_2;
  wire       [252:0]  mdsMatrix_7_3;
  wire       [253:0]  mdsMatrix_7_4;
  wire       [254:0]  mdsMatrix_7_5;
  wire       [252:0]  mdsMatrix_7_6;
  wire       [250:0]  mdsMatrix_7_7;
  wire       [253:0]  mdsMatrix_7_8;
  wire       [253:0]  mdsMatrix_8_0;
  wire       [254:0]  mdsMatrix_8_1;
  wire       [252:0]  mdsMatrix_8_2;
  wire       [253:0]  mdsMatrix_8_3;
  wire       [254:0]  mdsMatrix_8_4;
  wire       [252:0]  mdsMatrix_8_5;
  wire       [250:0]  mdsMatrix_8_6;
  wire       [253:0]  mdsMatrix_8_7;
  wire       [252:0]  mdsMatrix_8_8;
  wire       [3:0]    tempAddrVec_0;
  wire       [3:0]    tempAddrVec_1;
  wire       [3:0]    tempAddrVec_2;
  wire       [3:0]    tempAddrVec_3;
  wire       [3:0]    tempAddrVec_4;
  wire       [3:0]    tempAddrVec_5;
  wire       [3:0]    tempAddrVec_6;
  wire       [3:0]    tempAddrVec_7;
  wire       [3:0]    tempAddrVec_8;
  reg        [3:0]    io_addr_regNext;
  reg        [3:0]    io_addr_regNext_1;
  reg        [3:0]    io_addr_regNext_2;
  reg        [3:0]    io_addr_regNext_3;
  reg        [3:0]    io_addr_regNext_4;
  reg        [3:0]    io_addr_regNext_5;
  reg        [3:0]    io_addr_regNext_6;
  reg        [3:0]    io_addr_regNext_7;
  reg        [3:0]    io_addr_regNext_8;
  reg [254:0] mdsMem_0 [0:8];
  reg [254:0] mdsMem_1 [0:8];
  reg [254:0] mdsMem_2 [0:8];
  reg [254:0] mdsMem_3 [0:8];
  reg [254:0] mdsMem_4 [0:8];
  reg [254:0] mdsMem_5 [0:8];
  reg [254:0] mdsMem_6 [0:8];
  reg [254:0] mdsMem_7 [0:8];
  reg [254:0] mdsMem_8 [0:8];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  assign _zz_io_data_5 = 1'b1;
  assign _zz_io_data_6 = 1'b1;
  assign _zz_io_data_7 = 1'b1;
  assign _zz_io_data_8 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_16_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_16_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_16_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_16_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_16_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_16_mdsMem_5.bin",mdsMem_5);
  end
  always @(posedge clk) begin
    if(_zz_io_data_5) begin
      _zz_mdsMem_5_port0 <= mdsMem_5[tempAddrVec_5];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_16_mdsMem_6.bin",mdsMem_6);
  end
  always @(posedge clk) begin
    if(_zz_io_data_6) begin
      _zz_mdsMem_6_port0 <= mdsMem_6[tempAddrVec_6];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_16_mdsMem_7.bin",mdsMem_7);
  end
  always @(posedge clk) begin
    if(_zz_io_data_7) begin
      _zz_mdsMem_7_port0 <= mdsMem_7[tempAddrVec_7];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_16_mdsMem_8.bin",mdsMem_8);
  end
  always @(posedge clk) begin
    if(_zz_io_data_8) begin
      _zz_mdsMem_8_port0 <= mdsMem_8[tempAddrVec_8];
    end
  end

  assign mdsMatrix_0_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_0_1 = 250'h26a11bc2ae0808b28f46e64cadfa19888da1265cccd20cd0000000033333333;
  assign mdsMatrix_0_2 = 254'h2c59c154f04b2e0d209627474791ca2f8396d8008ba29c5ce8ba2e8b745d1746;
  assign mdsMatrix_0_3 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_0_4 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_0_5 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_0_6 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_0_7 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_0_8 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_1_0 = 250'h26a11bc2ae0808b28f46e64cadfa19888da1265cccd20cd0000000033333333;
  assign mdsMatrix_1_1 = 254'h2c59c154f04b2e0d209627474791ca2f8396d8008ba29c5ce8ba2e8b745d1746;
  assign mdsMatrix_1_2 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_1_3 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_1_4 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_1_5 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_1_6 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_1_7 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_1_8 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_2_0 = 254'h2c59c154f04b2e0d209627474791ca2f8396d8008ba29c5ce8ba2e8b745d1746;
  assign mdsMatrix_2_1 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_2_2 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_2_3 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_2_4 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_2_5 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_2_6 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_2_7 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_2_8 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_3_0 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_3_1 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_3_2 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_3_3 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_3_4 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_3_5 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_3_6 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_3_7 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_3_8 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_4_0 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign mdsMatrix_4_1 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_4_2 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_4_3 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_4_4 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_4_5 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_4_6 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_4_7 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_4_8 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_5_0 = 254'h336878f3307623cb7c59ab7002c086dcf35ac1256db6636d6db6db6d6db6db6e;
  assign mdsMatrix_5_1 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_5_2 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_5_3 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_5_4 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_5_5 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_5_6 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_5_7 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_5_8 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_6_0 = 255'h4ee5260a3853fe8ce81ed99de300fbbe930fcef08887a887ffffffff77777778;
  assign mdsMatrix_6_1 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_6_2 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_6_3 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_6_4 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_6_5 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_6_6 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_6_7 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_6_8 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_7_0 = 253'h1000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_7_1 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_7_2 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_7_3 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_7_4 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_7_5 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_7_6 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_7_7 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_7_8 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_8_0 = 254'h2a560940be7f68c5b1b341e3c607f697d777ea5b0f0eac3bffffffffc3c3c3c4;
  assign mdsMatrix_8_1 = 255'h686382243ccfd33827d7a80640616f2096770dc971c5d5c6555555548e38e38f;
  assign mdsMatrix_8_2 = 253'h1fc7355df918dde2fa9d580144e3a8d86b89bb94af2829791af286bc79435e51;
  assign mdsMatrix_8_3 = 254'h3b2bdc87aa3efee9ae1723366a40bcceee4bdb346665be65ffffffff9999999a;
  assign mdsMatrix_8_4 = 255'h48ea33132e2dec4a63f9ba4d5a60f73fbe266219f3ce60f3492492489e79e79f;
  assign mdsMatrix_8_5 = 253'h162ce0aa78259706904b13a3a3c8e517c1cb6c0045d14e2e745d1745ba2e8ba3;
  assign mdsMatrix_8_6 = 251'h6170efc625d5398afdc17ffa689a8b1daf7c1378590c4591642c8591642c859;
  assign mdsMatrix_8_7 = 254'h314f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_8_8 = 253'h1826c228b312e612e76d575d1fe038a47ab05b5c851e85eb6666666647ae147b;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign tempAddrVec_5 = io_addr_regNext_5;
  assign tempAddrVec_6 = io_addr_regNext_6;
  assign tempAddrVec_7 = io_addr_regNext_7;
  assign tempAddrVec_8 = io_addr_regNext_8;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  assign io_data_5 = _zz_mdsMem_5_port0;
  assign io_data_6 = _zz_mdsMem_6_port0;
  assign io_data_7 = _zz_mdsMem_7_port0;
  assign io_data_8 = _zz_mdsMem_8_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
    io_addr_regNext_5 <= io_addr;
    io_addr_regNext_6 <= io_addr;
    io_addr_regNext_7 <= io_addr;
    io_addr_regNext_8 <= io_addr;
  end


endmodule

module MatrixConstantMem_1 (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  output     [254:0]  io_data_3,
  output     [254:0]  io_data_4,
  input      [2:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  reg        [254:0]  _zz_mdsMem_3_port0;
  reg        [254:0]  _zz_mdsMem_4_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire                _zz_mdsMem_3_port;
  wire                _zz_io_data_3;
  wire                _zz_mdsMem_4_port;
  wire                _zz_io_data_4;
  wire       [250:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [254:0]  mdsMatrix_0_2;
  wire       [253:0]  mdsMatrix_0_3;
  wire       [254:0]  mdsMatrix_0_4;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [254:0]  mdsMatrix_1_1;
  wire       [253:0]  mdsMatrix_1_2;
  wire       [254:0]  mdsMatrix_1_3;
  wire       [249:0]  mdsMatrix_1_4;
  wire       [254:0]  mdsMatrix_2_0;
  wire       [253:0]  mdsMatrix_2_1;
  wire       [254:0]  mdsMatrix_2_2;
  wire       [249:0]  mdsMatrix_2_3;
  wire       [253:0]  mdsMatrix_2_4;
  wire       [253:0]  mdsMatrix_3_0;
  wire       [254:0]  mdsMatrix_3_1;
  wire       [249:0]  mdsMatrix_3_2;
  wire       [253:0]  mdsMatrix_3_3;
  wire       [254:0]  mdsMatrix_3_4;
  wire       [254:0]  mdsMatrix_4_0;
  wire       [249:0]  mdsMatrix_4_1;
  wire       [253:0]  mdsMatrix_4_2;
  wire       [254:0]  mdsMatrix_4_3;
  wire       [254:0]  mdsMatrix_4_4;
  wire       [2:0]    tempAddrVec_0;
  wire       [2:0]    tempAddrVec_1;
  wire       [2:0]    tempAddrVec_2;
  wire       [2:0]    tempAddrVec_3;
  wire       [2:0]    tempAddrVec_4;
  reg        [2:0]    io_addr_regNext;
  reg        [2:0]    io_addr_regNext_1;
  reg        [2:0]    io_addr_regNext_2;
  reg        [2:0]    io_addr_regNext_3;
  reg        [2:0]    io_addr_regNext_4;
  reg [254:0] mdsMem_0 [0:4];
  reg [254:0] mdsMem_1 [0:4];
  reg [254:0] mdsMem_2 [0:4];
  reg [254:0] mdsMem_3 [0:4];
  reg [254:0] mdsMem_4 [0:4];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  assign _zz_io_data_3 = 1'b1;
  assign _zz_io_data_4 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_15_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_15_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_15_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_15_mdsMem_3.bin",mdsMem_3);
  end
  always @(posedge clk) begin
    if(_zz_io_data_3) begin
      _zz_mdsMem_3_port0 <= mdsMem_3[tempAddrVec_3];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_15_mdsMem_4.bin",mdsMem_4);
  end
  always @(posedge clk) begin
    if(_zz_io_data_4) begin
      _zz_mdsMem_4_port0 <= mdsMem_4[tempAddrVec_4];
    end
  end

  assign mdsMatrix_0_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_0_1 = 255'h514f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_0_2 = 255'h66d0f1e660ec4796f8b356e005810db9e6b5824adb6cc6dadb6db6dadb6db6dc;
  assign mdsMatrix_0_3 = 254'h2000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_0_4 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_1_0 = 255'h514f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_1_1 = 255'h66d0f1e660ec4796f8b356e005810db9e6b5824adb6cc6dadb6db6dadb6db6dc;
  assign mdsMatrix_1_2 = 254'h2000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_1_3 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_1_4 = 250'h26a11bc2ae0808b28f46e64cadfa19888da1265cccd20cd0000000033333333;
  assign mdsMatrix_2_0 = 255'h66d0f1e660ec4796f8b356e005810db9e6b5824adb6cc6dadb6db6dadb6db6dc;
  assign mdsMatrix_2_1 = 254'h2000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_2_2 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_2_3 = 250'h26a11bc2ae0808b28f46e64cadfa19888da1265cccd20cd0000000033333333;
  assign mdsMatrix_2_4 = 254'h2c59c154f04b2e0d209627474791ca2f8396d8008ba29c5ce8ba2e8b745d1746;
  assign mdsMatrix_3_0 = 254'h2000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_3_1 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_3_2 = 250'h26a11bc2ae0808b28f46e64cadfa19888da1265cccd20cd0000000033333333;
  assign mdsMatrix_3_3 = 254'h2c59c154f04b2e0d209627474791ca2f8396d8008ba29c5ce8ba2e8b745d1746;
  assign mdsMatrix_3_4 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_4_0 = 255'h5cd95cf5500229281c7578047721063bd930778fe38d4f8daaaaaaaa1c71c71d;
  assign mdsMatrix_4_1 = 250'h26a11bc2ae0808b28f46e64cadfa19888da1265cccd20cd0000000033333333;
  assign mdsMatrix_4_2 = 254'h2c59c154f04b2e0d209627474791ca2f8396d8008ba29c5ce8ba2e8b745d1746;
  assign mdsMatrix_4_3 = 255'h629e6f8cc668fe30222690055bc13aae37d3c2acaaa992a9ffffffff55555556;
  assign mdsMatrix_4_4 = 255'h521d817b8c8fe0ff7e0b745318e0fe2a40c8936413b058ebc4ec4ec462762763;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign tempAddrVec_3 = io_addr_regNext_3;
  assign tempAddrVec_4 = io_addr_regNext_4;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  assign io_data_3 = _zz_mdsMem_3_port0;
  assign io_data_4 = _zz_mdsMem_4_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
    io_addr_regNext_3 <= io_addr;
    io_addr_regNext_4 <= io_addr;
  end


endmodule

module MatrixConstantMem (
  output     [254:0]  io_data_0,
  output     [254:0]  io_data_1,
  output     [254:0]  io_data_2,
  input      [1:0]    io_addr,
  input               clk,
  input               resetn
);

  reg        [254:0]  _zz_mdsMem_0_port0;
  reg        [254:0]  _zz_mdsMem_1_port0;
  reg        [254:0]  _zz_mdsMem_2_port0;
  wire                _zz_mdsMem_0_port;
  wire                _zz_io_data_0;
  wire                _zz_mdsMem_1_port;
  wire                _zz_io_data_1;
  wire                _zz_mdsMem_2_port;
  wire                _zz_io_data_2;
  wire       [253:0]  mdsMatrix_0_0;
  wire       [254:0]  mdsMatrix_0_1;
  wire       [250:0]  mdsMatrix_0_2;
  wire       [254:0]  mdsMatrix_1_0;
  wire       [250:0]  mdsMatrix_1_1;
  wire       [254:0]  mdsMatrix_1_2;
  wire       [250:0]  mdsMatrix_2_0;
  wire       [254:0]  mdsMatrix_2_1;
  wire       [254:0]  mdsMatrix_2_2;
  wire       [1:0]    tempAddrVec_0;
  wire       [1:0]    tempAddrVec_1;
  wire       [1:0]    tempAddrVec_2;
  reg        [1:0]    io_addr_regNext;
  reg        [1:0]    io_addr_regNext_1;
  reg        [1:0]    io_addr_regNext_2;
  reg [254:0] mdsMem_0 [0:2];
  reg [254:0] mdsMem_1 [0:2];
  reg [254:0] mdsMem_2 [0:2];

  assign _zz_io_data_0 = 1'b1;
  assign _zz_io_data_1 = 1'b1;
  assign _zz_io_data_2 = 1'b1;
  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_14_mdsMem_0.bin",mdsMem_0);
  end
  always @(posedge clk) begin
    if(_zz_io_data_0) begin
      _zz_mdsMem_0_port0 <= mdsMem_0[tempAddrVec_0];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_14_mdsMem_1.bin",mdsMem_1);
  end
  always @(posedge clk) begin
    if(_zz_io_data_1) begin
      _zz_mdsMem_1_port0 <= mdsMem_1[tempAddrVec_1];
    end
  end

  initial begin
    $readmemb("PoseidonTopLevel.v_toplevel_poseidonLoop_1_poseidonThread_1_mDSMatrixMultiplier_1_constants_matrixConstantMem_14_mdsMem_2.bin",mdsMem_2);
  end
  always @(posedge clk) begin
    if(_zz_io_data_2) begin
      _zz_mdsMem_2_port0 <= mdsMem_2[tempAddrVec_2];
    end
  end

  assign mdsMatrix_0_0 = 254'h2eb0c8399ccb80e7eeecb7fd521f62a8e4161ea9aaab36ab0000000055555555;
  assign mdsMatrix_0_1 = 255'h4000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_0_2 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_1_0 = 255'h4000000000000000000000000000000000000000000000000000000000000000;
  assign mdsMatrix_1_1 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_1_2 = 255'h514f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_2_0 = 251'h4d4237855c1011651e8dcc995bf433111b424cb999a419a0000000066666666;
  assign mdsMatrix_2_1 = 255'h514f37c663347f1811134802ade09d571be9e1565554c954ffffffffaaaaaaab;
  assign mdsMatrix_2_2 = 255'h66d0f1e660ec4796f8b356e005810db9e6b5824adb6cc6dadb6db6dadb6db6dc;
  assign tempAddrVec_0 = io_addr_regNext;
  assign tempAddrVec_1 = io_addr_regNext_1;
  assign tempAddrVec_2 = io_addr_regNext_2;
  assign io_data_0 = _zz_mdsMem_0_port0;
  assign io_data_1 = _zz_mdsMem_1_port0;
  assign io_data_2 = _zz_mdsMem_2_port0;
  always @(posedge clk) begin
    io_addr_regNext <= io_addr;
    io_addr_regNext_1 <= io_addr;
    io_addr_regNext_2 <= io_addr;
  end


endmodule

//SimAdderIP_22 replaced by SimAdderIP_22

module SimAdderIP_22 (
  input      [254:0]  io_inputA,
  input      [254:0]  io_inputB,
  output     [255:0]  io_outputS,
  input               clk,
  input               resetn
);

  wire       [255:0]  adderRes;
  wire       [255:0]  stages_0;
  reg        [255:0]  stages_1;
  reg        [255:0]  stages_2;
  reg        [255:0]  stages_3;
  reg        [255:0]  stages_4;
  reg        [255:0]  stages_5;
  reg        [255:0]  stages_6;
  reg        [255:0]  stages_7;
  reg        [255:0]  stages_8;
  reg        [255:0]  stages_9;
  reg        [255:0]  stages_10;
  reg        [255:0]  stages_11;
  reg        [255:0]  stages_12;
  reg        [255:0]  stages_13;
  reg        [255:0]  stages_14;
  reg        [255:0]  stages_15;
  reg        [255:0]  stages_16;

  assign adderRes = ({1'b0,io_inputA} + {1'b0,io_inputB});
  assign stages_0 = adderRes;
  assign io_outputS = stages_16;
  always @(posedge clk) begin
    stages_1 <= stages_0;
    stages_2 <= stages_1;
    stages_3 <= stages_2;
    stages_4 <= stages_3;
    stages_5 <= stages_4;
    stages_6 <= stages_5;
    stages_7 <= stages_6;
    stages_8 <= stages_7;
    stages_9 <= stages_8;
    stages_10 <= stages_9;
    stages_11 <= stages_10;
    stages_12 <= stages_11;
    stages_13 <= stages_12;
    stages_14 <= stages_13;
    stages_15 <= stages_14;
    stages_16 <= stages_15;
  end


endmodule

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

//SimAdderIP replaced by SimAdderIP

module SimAdderIP (
  input      [254:0]  io_inputA,
  input      [254:0]  io_inputB,
  output     [255:0]  io_outputS,
  input               clk,
  input               resetn
);

  wire       [255:0]  adderRes;
  wire       [255:0]  stages_0;
  reg        [255:0]  stages_1;
  reg        [255:0]  stages_2;
  reg        [255:0]  stages_3;
  reg        [255:0]  stages_4;
  reg        [255:0]  stages_5;
  reg        [255:0]  stages_6;
  reg        [255:0]  stages_7;
  reg        [255:0]  stages_8;

  assign adderRes = ({1'b0,io_inputA} + {1'b0,io_inputB});
  assign stages_0 = adderRes;
  assign io_outputS = stages_8;
  always @(posedge clk) begin
    stages_1 <= stages_0;
    stages_2 <= stages_1;
    stages_3 <= stages_2;
    stages_4 <= stages_3;
    stages_5 <= stages_4;
    stages_6 <= stages_5;
    stages_7 <= stages_6;
    stages_8 <= stages_7;
  end


endmodule

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

//MultiplierIPFlow replaced by MultiplierIPFlow

module MultiplierIPFlow (
  input               io_input_valid,
  input      [33:0]   io_input_payload_op1,
  input      [33:0]   io_input_payload_op2,
  output              io_output_valid,
  output     [67:0]   io_output_payload_res,
  input               clk,
  input               resetn
);

  wire       [67:0]   simMultiplierIP_1215_io_outputP;
  reg                 io_input_valid_delay_1;
  reg                 io_input_valid_delay_2;
  reg                 io_input_valid_delay_3;
  reg                 io_input_valid_delay_4;
  reg                 io_input_valid_delay_5;
  reg                 validPipe;

  SimMultiplierIP simMultiplierIP_1215 (
    .io_inputA     (io_input_payload_op1[33:0]             ), //i
    .io_inputB     (io_input_payload_op2[33:0]             ), //i
    .io_outputP    (simMultiplierIP_1215_io_outputP[67:0]  ), //o
    .clk           (clk                                    ), //i
    .resetn        (resetn                                 )  //i
  );
  assign io_output_valid = validPipe;
  assign io_output_payload_res = simMultiplierIP_1215_io_outputP;
  always @(posedge clk) begin
    if(!resetn) begin
      io_input_valid_delay_1 <= 1'b1;
      io_input_valid_delay_2 <= 1'b1;
      io_input_valid_delay_3 <= 1'b1;
      io_input_valid_delay_4 <= 1'b1;
      io_input_valid_delay_5 <= 1'b1;
      validPipe <= 1'b1;
    end else begin
      io_input_valid_delay_1 <= io_input_valid;
      io_input_valid_delay_2 <= io_input_valid_delay_1;
      io_input_valid_delay_3 <= io_input_valid_delay_2;
      io_input_valid_delay_4 <= io_input_valid_delay_3;
      io_input_valid_delay_5 <= io_input_valid_delay_4;
      validPipe <= io_input_valid_delay_5;
    end
  end


endmodule

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

//SimMultiplierIP replaced by SimMultiplierIP

module SimMultiplierIP (
  input      [33:0]   io_inputA,
  input      [33:0]   io_inputB,
  output     [67:0]   io_outputP,
  input               clk,
  input               resetn
);

  wire       [67:0]   _zz_mulRes;
  wire       [67:0]   mulRes;
  wire       [67:0]   stages_0;
  reg        [67:0]   stages_1;
  reg        [67:0]   stages_2;
  reg        [67:0]   stages_3;
  reg        [67:0]   stages_4;
  reg        [67:0]   stages_5;
  reg        [67:0]   stages_6;

  assign _zz_mulRes = (io_inputA * io_inputB);
  assign mulRes = _zz_mulRes;
  assign stages_0 = mulRes;
  assign io_outputP = stages_6;
  always @(posedge clk) begin
    stages_1 <= stages_0;
    stages_2 <= stages_1;
    stages_3 <= stages_2;
    stages_4 <= stages_3;
    stages_5 <= stages_4;
    stages_6 <= stages_5;
  end


endmodule
